module game_bar_rom
	(
		input wire clk,
		input wire [9:0] xpos,
		input wire [9:0] ypos,
		output reg [2:0] red,
		output reg [2:0] green,
		output reg [1:0] blue
	);

	(* rom_style = "block" *)


	reg [9:0] ypos_reg;
	reg [9:0] xpos_reg;

	always @(posedge clk)
		begin
		ypos_reg <= ypos;
		xpos_reg <= xpos;
		end

	always @*
	case ({xpos_reg, ypos_reg})
		20'b00011010100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011100110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011100110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011100110000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011101000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011101110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011110010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00011111110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100000010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100000010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100000100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100000100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100000110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100001000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100001010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100010000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100010000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100010000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100010000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100010000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100011010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100011010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100011010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100011010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100100000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100100000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100100000000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100100100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100100100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100100110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100101000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100101000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100101000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100110000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100110010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100110010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100110110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100110110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100110110000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100110110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100110110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b00100111000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000000000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000000000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000000010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000100000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000000100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000000100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000000100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000000110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001100000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000001100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000001110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000001110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000001110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000010010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000010010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000010010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000010010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000010010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000010010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000010100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000010110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000011000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000011010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000011100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000011100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000011110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000011110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000011110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100100000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000100110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000101010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000101010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000101010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000101010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000101100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000101100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000101100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000101110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000110010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000110010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000110100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000110110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000110110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000110110000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000110110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000110110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000111000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10000111000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111100000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10000111110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001000010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001000100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001000100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001000100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001000110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000110000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001000110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001001000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001001000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001001000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001001000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001001110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001001110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001010010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001010010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001010010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001010010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001010010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001010010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010100000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001010110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001010110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011100000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001011110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001011110000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001011110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001100010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001100100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001101000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101100000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101100000001010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001101100000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001101100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101100000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001101100000001111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001101100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001101100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001101110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110000000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110000000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110010000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110010000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110100000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110100000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110100000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110100000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110110000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110110000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110110000001011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001110110000001100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001110110000001101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001110110000001110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001110110000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001110110000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111000000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111000000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111000000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111010000001000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111010000001001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b10001111100000010000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001111100000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001111100000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		20'b10001111100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b00; end
		default: begin red <= 3'b000; green <= 3'b000; blue <= 2'b00; end
	endcase
endmodule