module pong_logo_rom
	(
		input wire clk,
		input wire [9:0] row,
		input wire [9:0] col,
		output reg [7:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [9:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		20'b00000011100000110100: color_data = 8'b10010010;
		20'b00000011100000110101: color_data = 8'b11011011;
		20'b00000011100000110110: color_data = 8'b11011011;
		20'b00000011100000110111: color_data = 8'b11011011;
		20'b00000011100000111000: color_data = 8'b11011011;
		20'b00000011100000111001: color_data = 8'b11011011;
		20'b00000011100000111010: color_data = 8'b11011011;
		20'b00000011100000111011: color_data = 8'b11011011;
		20'b00000011100000111100: color_data = 8'b11011011;
		20'b00000011100000111101: color_data = 8'b11011011;
		20'b00000011100000111110: color_data = 8'b11011011;
		20'b00000011100000111111: color_data = 8'b11011011;
		20'b00000011100001000000: color_data = 8'b11011011;
		20'b00000011100001000001: color_data = 8'b11011011;
		20'b00000011100001000010: color_data = 8'b11011011;
		20'b00000011100001000011: color_data = 8'b11011011;
		20'b00000011100001000100: color_data = 8'b11011011;
		20'b00000011100001000101: color_data = 8'b11011011;
		20'b00000011100001000110: color_data = 8'b11011011;
		20'b00000011100001000111: color_data = 8'b11011011;
		20'b00000011100001001000: color_data = 8'b11011011;
		20'b00000011100001001001: color_data = 8'b11011011;
		20'b00000011100001001010: color_data = 8'b11011011;
		20'b00000011100001001011: color_data = 8'b11011011;
		20'b00000011100001001100: color_data = 8'b11011011;
		20'b00000011100001001101: color_data = 8'b11011011;
		20'b00000011100001001110: color_data = 8'b11011011;
		20'b00000011100001001111: color_data = 8'b11011011;
		20'b00000011100001010000: color_data = 8'b11011011;
		20'b00000011100001010001: color_data = 8'b11011011;
		20'b00000011100001010010: color_data = 8'b11011011;
		20'b00000011100001010011: color_data = 8'b11011011;
		20'b00000011100001010100: color_data = 8'b11011011;
		20'b00000011100001010101: color_data = 8'b11011011;
		20'b00000011100001010110: color_data = 8'b11011011;
		20'b00000011100001010111: color_data = 8'b11011011;
		20'b00000011100001011000: color_data = 8'b11011011;
		20'b00000011100001011001: color_data = 8'b11011011;
		20'b00000011100001011010: color_data = 8'b11011011;
		20'b00000011100001011011: color_data = 8'b11011011;
		20'b00000011100001011100: color_data = 8'b11011011;
		20'b00000011100001011101: color_data = 8'b11011011;
		20'b00000011100001011110: color_data = 8'b11011011;
		20'b00000011100001011111: color_data = 8'b11011011;
		20'b00000011100001100000: color_data = 8'b11011011;
		20'b00000011100001100001: color_data = 8'b11011011;
		20'b00000011100001100010: color_data = 8'b11011011;
		20'b00000011100001100011: color_data = 8'b11011011;

		20'b00000011110000110100: color_data = 8'b11011011;
		20'b00000011110000110101: color_data = 8'b11111111;
		20'b00000011110000110110: color_data = 8'b11111111;
		20'b00000011110000110111: color_data = 8'b11111111;
		20'b00000011110000111000: color_data = 8'b11111111;
		20'b00000011110000111001: color_data = 8'b11111111;
		20'b00000011110000111010: color_data = 8'b11111111;
		20'b00000011110000111011: color_data = 8'b11111111;
		20'b00000011110000111100: color_data = 8'b11111111;
		20'b00000011110000111101: color_data = 8'b11111111;
		20'b00000011110000111110: color_data = 8'b11111111;
		20'b00000011110000111111: color_data = 8'b11111111;
		20'b00000011110001000000: color_data = 8'b11111111;
		20'b00000011110001000001: color_data = 8'b11111111;
		20'b00000011110001000010: color_data = 8'b11111111;
		20'b00000011110001000011: color_data = 8'b11111111;
		20'b00000011110001000100: color_data = 8'b11111111;
		20'b00000011110001000101: color_data = 8'b11111111;
		20'b00000011110001000110: color_data = 8'b11111111;
		20'b00000011110001000111: color_data = 8'b11111111;
		20'b00000011110001001000: color_data = 8'b11111111;
		20'b00000011110001001001: color_data = 8'b11111111;
		20'b00000011110001001010: color_data = 8'b11111111;
		20'b00000011110001001011: color_data = 8'b11111111;
		20'b00000011110001001100: color_data = 8'b11111111;
		20'b00000011110001001101: color_data = 8'b11111111;
		20'b00000011110001001110: color_data = 8'b11111111;
		20'b00000011110001001111: color_data = 8'b11111111;
		20'b00000011110001010000: color_data = 8'b11111111;
		20'b00000011110001010001: color_data = 8'b11111111;
		20'b00000011110001010010: color_data = 8'b11111111;
		20'b00000011110001010011: color_data = 8'b11111111;
		20'b00000011110001010100: color_data = 8'b11111111;
		20'b00000011110001010101: color_data = 8'b11111111;
		20'b00000011110001010110: color_data = 8'b11111111;
		20'b00000011110001010111: color_data = 8'b11111111;
		20'b00000011110001011000: color_data = 8'b11111111;
		20'b00000011110001011001: color_data = 8'b11111111;
		20'b00000011110001011010: color_data = 8'b11111111;
		20'b00000011110001011011: color_data = 8'b11111111;
		20'b00000011110001011100: color_data = 8'b11111111;
		20'b00000011110001011101: color_data = 8'b11111111;
		20'b00000011110001011110: color_data = 8'b11111111;
		20'b00000011110001011111: color_data = 8'b11111111;
		20'b00000011110001100000: color_data = 8'b11111111;
		20'b00000011110001100001: color_data = 8'b11111111;
		20'b00000011110001100010: color_data = 8'b11111111;
		20'b00000011110001100011: color_data = 8'b11111111;

		20'b00000100000000110100: color_data = 8'b11011011;
		20'b00000100000000110101: color_data = 8'b11111111;
		20'b00000100000000110110: color_data = 8'b11111111;
		20'b00000100000000110111: color_data = 8'b11111111;
		20'b00000100000000111000: color_data = 8'b11111111;
		20'b00000100000000111001: color_data = 8'b11111111;
		20'b00000100000000111010: color_data = 8'b11111111;
		20'b00000100000000111011: color_data = 8'b11111111;
		20'b00000100000000111100: color_data = 8'b11111111;
		20'b00000100000000111101: color_data = 8'b11111111;
		20'b00000100000000111110: color_data = 8'b11111111;
		20'b00000100000000111111: color_data = 8'b11111111;
		20'b00000100000001000000: color_data = 8'b11111111;
		20'b00000100000001000001: color_data = 8'b11111111;
		20'b00000100000001000010: color_data = 8'b11111111;
		20'b00000100000001000011: color_data = 8'b11111111;
		20'b00000100000001000100: color_data = 8'b11111111;
		20'b00000100000001000101: color_data = 8'b11111111;
		20'b00000100000001000110: color_data = 8'b11111111;
		20'b00000100000001000111: color_data = 8'b11111111;
		20'b00000100000001001000: color_data = 8'b11111111;
		20'b00000100000001001001: color_data = 8'b11111111;
		20'b00000100000001001010: color_data = 8'b11111111;
		20'b00000100000001001011: color_data = 8'b11111111;
		20'b00000100000001001100: color_data = 8'b11111111;
		20'b00000100000001001101: color_data = 8'b11111111;
		20'b00000100000001001110: color_data = 8'b11111111;
		20'b00000100000001001111: color_data = 8'b11111111;
		20'b00000100000001010000: color_data = 8'b11111111;
		20'b00000100000001010001: color_data = 8'b11111111;
		20'b00000100000001010010: color_data = 8'b11111111;
		20'b00000100000001010011: color_data = 8'b11111111;
		20'b00000100000001010100: color_data = 8'b11111111;
		20'b00000100000001010101: color_data = 8'b11111111;
		20'b00000100000001010110: color_data = 8'b11111111;
		20'b00000100000001010111: color_data = 8'b11111111;
		20'b00000100000001011000: color_data = 8'b11111111;
		20'b00000100000001011001: color_data = 8'b11111111;
		20'b00000100000001011010: color_data = 8'b11111111;
		20'b00000100000001011011: color_data = 8'b11111111;
		20'b00000100000001011100: color_data = 8'b11111111;
		20'b00000100000001011101: color_data = 8'b11111111;
		20'b00000100000001011110: color_data = 8'b11111111;
		20'b00000100000001011111: color_data = 8'b11111111;
		20'b00000100000001100000: color_data = 8'b11111111;
		20'b00000100000001100001: color_data = 8'b11111111;
		20'b00000100000001100010: color_data = 8'b11111111;
		20'b00000100000001100011: color_data = 8'b11111111;

		20'b00000100010000110100: color_data = 8'b11011011;
		20'b00000100010000110101: color_data = 8'b11111111;
		20'b00000100010000110110: color_data = 8'b11111111;
		20'b00000100010000110111: color_data = 8'b11111111;
		20'b00000100010000111000: color_data = 8'b11111111;
		20'b00000100010000111001: color_data = 8'b11111111;
		20'b00000100010000111010: color_data = 8'b11111111;
		20'b00000100010000111011: color_data = 8'b11111111;
		20'b00000100010000111100: color_data = 8'b11111111;
		20'b00000100010000111101: color_data = 8'b11111111;
		20'b00000100010000111110: color_data = 8'b11111111;
		20'b00000100010000111111: color_data = 8'b11111111;
		20'b00000100010001000000: color_data = 8'b11111111;
		20'b00000100010001000001: color_data = 8'b11111111;
		20'b00000100010001000010: color_data = 8'b11111111;
		20'b00000100010001000011: color_data = 8'b11111111;
		20'b00000100010001000100: color_data = 8'b11111111;
		20'b00000100010001000101: color_data = 8'b11111111;
		20'b00000100010001000110: color_data = 8'b11111111;
		20'b00000100010001000111: color_data = 8'b11111111;
		20'b00000100010001001000: color_data = 8'b11111111;
		20'b00000100010001001001: color_data = 8'b11111111;
		20'b00000100010001001010: color_data = 8'b11111111;
		20'b00000100010001001011: color_data = 8'b11111111;
		20'b00000100010001001100: color_data = 8'b11111111;
		20'b00000100010001001101: color_data = 8'b11111111;
		20'b00000100010001001110: color_data = 8'b11111111;
		20'b00000100010001001111: color_data = 8'b11111111;
		20'b00000100010001010000: color_data = 8'b11111111;
		20'b00000100010001010001: color_data = 8'b11111111;
		20'b00000100010001010010: color_data = 8'b11111111;
		20'b00000100010001010011: color_data = 8'b11111111;
		20'b00000100010001010100: color_data = 8'b11111111;
		20'b00000100010001010101: color_data = 8'b11111111;
		20'b00000100010001010110: color_data = 8'b11111111;
		20'b00000100010001010111: color_data = 8'b11111111;
		20'b00000100010001011000: color_data = 8'b11111111;
		20'b00000100010001011001: color_data = 8'b11111111;
		20'b00000100010001011010: color_data = 8'b11111111;
		20'b00000100010001011011: color_data = 8'b11111111;
		20'b00000100010001011100: color_data = 8'b11111111;
		20'b00000100010001011101: color_data = 8'b11111111;
		20'b00000100010001011110: color_data = 8'b11111111;
		20'b00000100010001011111: color_data = 8'b11111111;
		20'b00000100010001100000: color_data = 8'b11111111;
		20'b00000100010001100001: color_data = 8'b11111111;
		20'b00000100010001100010: color_data = 8'b11111111;
		20'b00000100010001100011: color_data = 8'b11111111;

		20'b00000100100000110100: color_data = 8'b11011011;
		20'b00000100100000110101: color_data = 8'b11111111;
		20'b00000100100000110110: color_data = 8'b11111111;
		20'b00000100100000110111: color_data = 8'b11111111;
		20'b00000100100000111000: color_data = 8'b11111111;
		20'b00000100100000111001: color_data = 8'b11111111;
		20'b00000100100000111010: color_data = 8'b11111111;
		20'b00000100100000111011: color_data = 8'b11111111;
		20'b00000100100000111100: color_data = 8'b11111111;
		20'b00000100100000111101: color_data = 8'b11111111;
		20'b00000100100000111110: color_data = 8'b11111111;
		20'b00000100100000111111: color_data = 8'b11111111;
		20'b00000100100001000000: color_data = 8'b11111111;
		20'b00000100100001000001: color_data = 8'b11111111;
		20'b00000100100001000010: color_data = 8'b11111111;
		20'b00000100100001000011: color_data = 8'b11111111;
		20'b00000100100001000100: color_data = 8'b11111111;
		20'b00000100100001000101: color_data = 8'b11111111;
		20'b00000100100001000110: color_data = 8'b11111111;
		20'b00000100100001000111: color_data = 8'b11111111;
		20'b00000100100001001000: color_data = 8'b11111111;
		20'b00000100100001001001: color_data = 8'b11111111;
		20'b00000100100001001010: color_data = 8'b11111111;
		20'b00000100100001001011: color_data = 8'b11111111;
		20'b00000100100001001100: color_data = 8'b11111111;
		20'b00000100100001001101: color_data = 8'b11111111;
		20'b00000100100001001110: color_data = 8'b11111111;
		20'b00000100100001001111: color_data = 8'b11111111;
		20'b00000100100001010000: color_data = 8'b11111111;
		20'b00000100100001010001: color_data = 8'b11111111;
		20'b00000100100001010010: color_data = 8'b11111111;
		20'b00000100100001010011: color_data = 8'b11111111;
		20'b00000100100001010100: color_data = 8'b11111111;
		20'b00000100100001010101: color_data = 8'b11111111;
		20'b00000100100001010110: color_data = 8'b11111111;
		20'b00000100100001010111: color_data = 8'b11111111;
		20'b00000100100001011000: color_data = 8'b11111111;
		20'b00000100100001011001: color_data = 8'b11111111;
		20'b00000100100001011010: color_data = 8'b11111111;
		20'b00000100100001011011: color_data = 8'b11111111;
		20'b00000100100001011100: color_data = 8'b11111111;
		20'b00000100100001011101: color_data = 8'b11111111;
		20'b00000100100001011110: color_data = 8'b11111111;
		20'b00000100100001011111: color_data = 8'b11111111;
		20'b00000100100001100000: color_data = 8'b11111111;
		20'b00000100100001100001: color_data = 8'b11111111;
		20'b00000100100001100010: color_data = 8'b11111111;
		20'b00000100100001100011: color_data = 8'b11111111;

		20'b00000100110000110100: color_data = 8'b11011011;
		20'b00000100110000110101: color_data = 8'b11111111;
		20'b00000100110000110110: color_data = 8'b11111111;
		20'b00000100110000110111: color_data = 8'b11111111;
		20'b00000100110000111000: color_data = 8'b11111111;
		20'b00000100110000111001: color_data = 8'b11111111;
		20'b00000100110000111010: color_data = 8'b11111111;
		20'b00000100110000111011: color_data = 8'b11111111;
		20'b00000100110000111100: color_data = 8'b11111111;
		20'b00000100110000111101: color_data = 8'b11111111;
		20'b00000100110000111110: color_data = 8'b11111111;
		20'b00000100110000111111: color_data = 8'b11111111;
		20'b00000100110001000000: color_data = 8'b11111111;
		20'b00000100110001000001: color_data = 8'b11111111;
		20'b00000100110001000010: color_data = 8'b11111111;
		20'b00000100110001000011: color_data = 8'b11111111;
		20'b00000100110001000100: color_data = 8'b11111111;
		20'b00000100110001000101: color_data = 8'b11111111;
		20'b00000100110001000110: color_data = 8'b11111111;
		20'b00000100110001000111: color_data = 8'b11111111;
		20'b00000100110001001000: color_data = 8'b11111111;
		20'b00000100110001001001: color_data = 8'b11111111;
		20'b00000100110001001010: color_data = 8'b11111111;
		20'b00000100110001001011: color_data = 8'b11111111;
		20'b00000100110001001100: color_data = 8'b11111111;
		20'b00000100110001001101: color_data = 8'b11111111;
		20'b00000100110001001110: color_data = 8'b11111111;
		20'b00000100110001001111: color_data = 8'b11111111;
		20'b00000100110001010000: color_data = 8'b11111111;
		20'b00000100110001010001: color_data = 8'b11111111;
		20'b00000100110001010010: color_data = 8'b11111111;
		20'b00000100110001010011: color_data = 8'b11111111;
		20'b00000100110001010100: color_data = 8'b11111111;
		20'b00000100110001010101: color_data = 8'b11111111;
		20'b00000100110001010110: color_data = 8'b11111111;
		20'b00000100110001010111: color_data = 8'b11111111;
		20'b00000100110001011000: color_data = 8'b11111111;
		20'b00000100110001011001: color_data = 8'b11111111;
		20'b00000100110001011010: color_data = 8'b11111111;
		20'b00000100110001011011: color_data = 8'b11111111;
		20'b00000100110001011100: color_data = 8'b11111111;
		20'b00000100110001011101: color_data = 8'b11111111;
		20'b00000100110001011110: color_data = 8'b11111111;
		20'b00000100110001011111: color_data = 8'b11111111;
		20'b00000100110001100000: color_data = 8'b11111111;
		20'b00000100110001100001: color_data = 8'b11111111;
		20'b00000100110001100010: color_data = 8'b11111111;
		20'b00000100110001100011: color_data = 8'b11111111;

		20'b00000101000000110100: color_data = 8'b11011011;
		20'b00000101000000110101: color_data = 8'b11111111;
		20'b00000101000000110110: color_data = 8'b11111111;
		20'b00000101000000110111: color_data = 8'b11111111;
		20'b00000101000000111000: color_data = 8'b11111111;
		20'b00000101000000111001: color_data = 8'b11111111;
		20'b00000101000000111010: color_data = 8'b11111111;
		20'b00000101000000111011: color_data = 8'b11111111;
		20'b00000101000000111100: color_data = 8'b11111111;
		20'b00000101000000111101: color_data = 8'b11111111;
		20'b00000101000000111110: color_data = 8'b11111111;
		20'b00000101000000111111: color_data = 8'b11111111;
		20'b00000101000001000000: color_data = 8'b11111111;
		20'b00000101000001000001: color_data = 8'b11111111;
		20'b00000101000001000010: color_data = 8'b11111111;
		20'b00000101000001000011: color_data = 8'b11111111;
		20'b00000101000001000100: color_data = 8'b11111111;
		20'b00000101000001000101: color_data = 8'b11111111;
		20'b00000101000001000110: color_data = 8'b11111111;
		20'b00000101000001000111: color_data = 8'b11111111;
		20'b00000101000001001000: color_data = 8'b11111111;
		20'b00000101000001001001: color_data = 8'b11111111;
		20'b00000101000001001010: color_data = 8'b11111111;
		20'b00000101000001001011: color_data = 8'b11111111;
		20'b00000101000001001100: color_data = 8'b11111111;
		20'b00000101000001001101: color_data = 8'b11111111;
		20'b00000101000001001110: color_data = 8'b11111111;
		20'b00000101000001001111: color_data = 8'b11111111;
		20'b00000101000001010000: color_data = 8'b11111111;
		20'b00000101000001010001: color_data = 8'b11111111;
		20'b00000101000001010010: color_data = 8'b11111111;
		20'b00000101000001010011: color_data = 8'b11111111;
		20'b00000101000001010100: color_data = 8'b11111111;
		20'b00000101000001010101: color_data = 8'b11111111;
		20'b00000101000001010110: color_data = 8'b11111111;
		20'b00000101000001010111: color_data = 8'b11111111;
		20'b00000101000001011000: color_data = 8'b11111111;
		20'b00000101000001011001: color_data = 8'b11111111;
		20'b00000101000001011010: color_data = 8'b11111111;
		20'b00000101000001011011: color_data = 8'b11111111;
		20'b00000101000001011100: color_data = 8'b11111111;
		20'b00000101000001011101: color_data = 8'b11111111;
		20'b00000101000001011110: color_data = 8'b11111111;
		20'b00000101000001011111: color_data = 8'b11111111;
		20'b00000101000001100000: color_data = 8'b11111111;
		20'b00000101000001100001: color_data = 8'b11111111;
		20'b00000101000001100010: color_data = 8'b11111111;
		20'b00000101000001100011: color_data = 8'b11111111;

		20'b00000101010000110100: color_data = 8'b11011011;
		20'b00000101010000110101: color_data = 8'b11111111;
		20'b00000101010000110110: color_data = 8'b11111111;
		20'b00000101010000110111: color_data = 8'b11111111;
		20'b00000101010000111000: color_data = 8'b11111111;
		20'b00000101010000111001: color_data = 8'b11111111;
		20'b00000101010000111010: color_data = 8'b11111111;
		20'b00000101010000111011: color_data = 8'b11111111;
		20'b00000101010000111100: color_data = 8'b11111111;
		20'b00000101010000111101: color_data = 8'b11111111;
		20'b00000101010000111110: color_data = 8'b11111111;
		20'b00000101010000111111: color_data = 8'b11111111;
		20'b00000101010001000000: color_data = 8'b11111111;
		20'b00000101010001000001: color_data = 8'b11111111;
		20'b00000101010001000010: color_data = 8'b11111111;
		20'b00000101010001000011: color_data = 8'b11111111;
		20'b00000101010001000100: color_data = 8'b11111111;
		20'b00000101010001000101: color_data = 8'b11111111;
		20'b00000101010001000110: color_data = 8'b11111111;
		20'b00000101010001000111: color_data = 8'b11111111;
		20'b00000101010001001000: color_data = 8'b11111111;
		20'b00000101010001001001: color_data = 8'b11111111;
		20'b00000101010001001010: color_data = 8'b11111111;
		20'b00000101010001001011: color_data = 8'b11111111;
		20'b00000101010001001100: color_data = 8'b11111111;
		20'b00000101010001001101: color_data = 8'b11111111;
		20'b00000101010001001110: color_data = 8'b11111111;
		20'b00000101010001001111: color_data = 8'b11111111;
		20'b00000101010001010000: color_data = 8'b11111111;
		20'b00000101010001010001: color_data = 8'b11111111;
		20'b00000101010001010010: color_data = 8'b11111111;
		20'b00000101010001010011: color_data = 8'b11111111;
		20'b00000101010001010100: color_data = 8'b11111111;
		20'b00000101010001010101: color_data = 8'b11111111;
		20'b00000101010001010110: color_data = 8'b11111111;
		20'b00000101010001010111: color_data = 8'b11111111;
		20'b00000101010001011000: color_data = 8'b11111111;
		20'b00000101010001011001: color_data = 8'b11111111;
		20'b00000101010001011010: color_data = 8'b11111111;
		20'b00000101010001011011: color_data = 8'b11111111;
		20'b00000101010001011100: color_data = 8'b11111111;
		20'b00000101010001011101: color_data = 8'b11111111;
		20'b00000101010001011110: color_data = 8'b11111111;
		20'b00000101010001011111: color_data = 8'b11111111;
		20'b00000101010001100000: color_data = 8'b11111111;
		20'b00000101010001100001: color_data = 8'b11111111;
		20'b00000101010001100010: color_data = 8'b11111111;
		20'b00000101010001100011: color_data = 8'b11111111;

		20'b00000101100000110100: color_data = 8'b11011011;
		20'b00000101100000110101: color_data = 8'b11111111;
		20'b00000101100000110110: color_data = 8'b11111111;
		20'b00000101100000110111: color_data = 8'b11111111;
		20'b00000101100000111000: color_data = 8'b11111111;
		20'b00000101100000111001: color_data = 8'b11111111;
		20'b00000101100000111010: color_data = 8'b11111111;
		20'b00000101100000111011: color_data = 8'b11111111;
		20'b00000101100000111100: color_data = 8'b11111111;
		20'b00000101100000111101: color_data = 8'b11111111;
		20'b00000101100000111110: color_data = 8'b11111111;
		20'b00000101100000111111: color_data = 8'b11111111;
		20'b00000101100001000000: color_data = 8'b11111111;
		20'b00000101100001000001: color_data = 8'b11111111;
		20'b00000101100001000010: color_data = 8'b11111111;
		20'b00000101100001000011: color_data = 8'b11111111;
		20'b00000101100001000100: color_data = 8'b11111111;
		20'b00000101100001000101: color_data = 8'b11111111;
		20'b00000101100001000110: color_data = 8'b11111111;
		20'b00000101100001000111: color_data = 8'b11111111;
		20'b00000101100001001000: color_data = 8'b11111111;
		20'b00000101100001001001: color_data = 8'b11111111;
		20'b00000101100001001010: color_data = 8'b11111111;
		20'b00000101100001001011: color_data = 8'b11111111;
		20'b00000101100001001100: color_data = 8'b11111111;
		20'b00000101100001001101: color_data = 8'b11111111;
		20'b00000101100001001110: color_data = 8'b11111111;
		20'b00000101100001001111: color_data = 8'b11111111;
		20'b00000101100001010000: color_data = 8'b11111111;
		20'b00000101100001010001: color_data = 8'b11111111;
		20'b00000101100001010010: color_data = 8'b11111111;
		20'b00000101100001010011: color_data = 8'b11111111;
		20'b00000101100001010100: color_data = 8'b11111111;
		20'b00000101100001010101: color_data = 8'b11111111;
		20'b00000101100001010110: color_data = 8'b11111111;
		20'b00000101100001010111: color_data = 8'b11111111;
		20'b00000101100001011000: color_data = 8'b11111111;
		20'b00000101100001011001: color_data = 8'b11111111;
		20'b00000101100001011010: color_data = 8'b11111111;
		20'b00000101100001011011: color_data = 8'b11111111;
		20'b00000101100001011100: color_data = 8'b11111111;
		20'b00000101100001011101: color_data = 8'b11111111;
		20'b00000101100001011110: color_data = 8'b11111111;
		20'b00000101100001011111: color_data = 8'b11111111;
		20'b00000101100001100000: color_data = 8'b11111111;
		20'b00000101100001100001: color_data = 8'b11111111;
		20'b00000101100001100010: color_data = 8'b11111111;
		20'b00000101100001100011: color_data = 8'b11111111;

		20'b00000101110000110100: color_data = 8'b11011011;
		20'b00000101110000110101: color_data = 8'b11011011;
		20'b00000101110000110110: color_data = 8'b11011011;
		20'b00000101110000110111: color_data = 8'b11011011;
		20'b00000101110000111000: color_data = 8'b11011011;
		20'b00000101110000111001: color_data = 8'b11011011;
		20'b00000101110000111010: color_data = 8'b11011011;
		20'b00000101110000111011: color_data = 8'b11011011;
		20'b00000101110000111100: color_data = 8'b11011011;
		20'b00000101110000111101: color_data = 8'b11011011;
		20'b00000101110000111110: color_data = 8'b11011011;
		20'b00000101110000111111: color_data = 8'b11011011;
		20'b00000101110001000000: color_data = 8'b11011011;
		20'b00000101110001000001: color_data = 8'b11011011;
		20'b00000101110001000010: color_data = 8'b11011011;
		20'b00000101110001000011: color_data = 8'b11011011;
		20'b00000101110001000100: color_data = 8'b11011011;
		20'b00000101110001000101: color_data = 8'b11011011;
		20'b00000101110001000110: color_data = 8'b11011011;
		20'b00000101110001000111: color_data = 8'b11011011;
		20'b00000101110001001000: color_data = 8'b11011011;
		20'b00000101110001001001: color_data = 8'b11011011;
		20'b00000101110001001010: color_data = 8'b11011011;
		20'b00000101110001001011: color_data = 8'b11011011;
		20'b00000101110001001100: color_data = 8'b11011011;
		20'b00000101110001001101: color_data = 8'b11011011;
		20'b00000101110001001110: color_data = 8'b11011011;
		20'b00000101110001001111: color_data = 8'b11011011;
		20'b00000101110001010000: color_data = 8'b11011011;
		20'b00000101110001010001: color_data = 8'b11011011;
		20'b00000101110001010010: color_data = 8'b11011011;
		20'b00000101110001010011: color_data = 8'b11011011;
		20'b00000101110001010100: color_data = 8'b11011011;
		20'b00000101110001010101: color_data = 8'b11011011;
		20'b00000101110001010110: color_data = 8'b11011011;
		20'b00000101110001010111: color_data = 8'b11011011;
		20'b00000101110001011000: color_data = 8'b11011011;
		20'b00000101110001011001: color_data = 8'b11011011;
		20'b00000101110001011010: color_data = 8'b11011011;
		20'b00000101110001011011: color_data = 8'b11011011;
		20'b00000101110001011100: color_data = 8'b11011011;
		20'b00000101110001011101: color_data = 8'b11011011;
		20'b00000101110001011110: color_data = 8'b11011011;
		20'b00000101110001011111: color_data = 8'b11011011;
		20'b00000101110001100000: color_data = 8'b11011011;
		20'b00000101110001100001: color_data = 8'b11011011;
		20'b00000101110001100010: color_data = 8'b11011011;
		20'b00000101110001100011: color_data = 8'b11111111;

		20'b00010011000000001001: color_data = 8'b11011011;
		20'b00010011000000001010: color_data = 8'b11011011;
		20'b00010011000000001011: color_data = 8'b11011011;
		20'b00010011000000001100: color_data = 8'b11011011;
		20'b00010011000000001101: color_data = 8'b11011011;
		20'b00010011000000001110: color_data = 8'b11011011;
		20'b00010011000000001111: color_data = 8'b11011011;
		20'b00010011000000010000: color_data = 8'b11011011;
		20'b00010011000000010001: color_data = 8'b11011011;
		20'b00010011000000010010: color_data = 8'b11011011;
		20'b00010011000000010011: color_data = 8'b11011011;
		20'b00010011000000010100: color_data = 8'b11011011;
		20'b00010011000000010101: color_data = 8'b11011011;
		20'b00010011000000010110: color_data = 8'b11011011;
		20'b00010011000000010111: color_data = 8'b11011011;
		20'b00010011000000011000: color_data = 8'b11011011;
		20'b00010011000000011001: color_data = 8'b11011011;
		20'b00010011000000011010: color_data = 8'b11011011;
		20'b00010011000000011011: color_data = 8'b11011011;
		20'b00010011000000011100: color_data = 8'b11011011;
		20'b00010011000000011101: color_data = 8'b11011011;
		20'b00010011000000011110: color_data = 8'b11011011;
		20'b00010011000000011111: color_data = 8'b11011011;
		20'b00010011000000100000: color_data = 8'b11011011;
		20'b00010011000000100001: color_data = 8'b11011011;
		20'b00010011000000100010: color_data = 8'b11011011;
		20'b00010011000000100011: color_data = 8'b11011011;
		20'b00010011000000100100: color_data = 8'b11011011;
		20'b00010011000000100101: color_data = 8'b11011011;
		20'b00010011000000100110: color_data = 8'b11011011;
		20'b00010011000000100111: color_data = 8'b11011011;
		20'b00010011000000101000: color_data = 8'b11011011;
		20'b00010011000000101001: color_data = 8'b11011011;
		20'b00010011000000101010: color_data = 8'b11011011;
		20'b00010011000000101011: color_data = 8'b11011011;
		20'b00010011000000101100: color_data = 8'b11011011;
		20'b00010011000000101101: color_data = 8'b11011011;
		20'b00010011000000101110: color_data = 8'b11011011;
		20'b00010011000000101111: color_data = 8'b11011011;
		20'b00010011000000111001: color_data = 8'b11011011;
		20'b00010011000000111010: color_data = 8'b11011011;
		20'b00010011000000111011: color_data = 8'b11011011;
		20'b00010011000000111100: color_data = 8'b11011011;
		20'b00010011000000111101: color_data = 8'b11011011;
		20'b00010011000000111110: color_data = 8'b11011011;
		20'b00010011000000111111: color_data = 8'b11011011;
		20'b00010011000001000000: color_data = 8'b11011011;
		20'b00010011000001000001: color_data = 8'b11011011;
		20'b00010011000001000010: color_data = 8'b11011011;
		20'b00010011000001000011: color_data = 8'b11011011;
		20'b00010011000001000100: color_data = 8'b11011011;
		20'b00010011000001000101: color_data = 8'b11011011;
		20'b00010011000001000110: color_data = 8'b11011011;
		20'b00010011000001000111: color_data = 8'b11011011;
		20'b00010011000001001000: color_data = 8'b11011011;
		20'b00010011000001001001: color_data = 8'b11011011;
		20'b00010011000001001010: color_data = 8'b11011011;
		20'b00010011000001001011: color_data = 8'b11011011;
		20'b00010011000001001100: color_data = 8'b11011011;
		20'b00010011000001001101: color_data = 8'b11011011;
		20'b00010011000001001110: color_data = 8'b11011011;
		20'b00010011000001001111: color_data = 8'b11011011;
		20'b00010011000001010000: color_data = 8'b11011011;
		20'b00010011000001010001: color_data = 8'b11011011;
		20'b00010011000001010010: color_data = 8'b11011011;
		20'b00010011000001010011: color_data = 8'b11011011;
		20'b00010011000001010100: color_data = 8'b11011011;
		20'b00010011000001010101: color_data = 8'b11011011;
		20'b00010011000001010110: color_data = 8'b11011011;
		20'b00010011000001010111: color_data = 8'b11011011;
		20'b00010011000001011000: color_data = 8'b11011011;
		20'b00010011000001011001: color_data = 8'b11011011;
		20'b00010011000001011010: color_data = 8'b11011011;
		20'b00010011000001011011: color_data = 8'b11011011;
		20'b00010011000001011100: color_data = 8'b11011011;
		20'b00010011000001011101: color_data = 8'b11011011;
		20'b00010011000001011110: color_data = 8'b11011011;
		20'b00010011000001011111: color_data = 8'b10010010;
		20'b00010011000001101000: color_data = 8'b10010010;
		20'b00010011000001101001: color_data = 8'b11011011;
		20'b00010011000001101010: color_data = 8'b11011011;
		20'b00010011000001101011: color_data = 8'b11011011;
		20'b00010011000001101100: color_data = 8'b11011011;
		20'b00010011000001101101: color_data = 8'b11011011;
		20'b00010011000001101110: color_data = 8'b11011011;
		20'b00010011000001101111: color_data = 8'b11011011;
		20'b00010011000001110000: color_data = 8'b11011011;
		20'b00010011000001110001: color_data = 8'b11011011;
		20'b00010011000001110010: color_data = 8'b11011011;
		20'b00010011000001110011: color_data = 8'b11011011;
		20'b00010011000001110100: color_data = 8'b11011011;
		20'b00010011000001110101: color_data = 8'b11011011;
		20'b00010011000001110110: color_data = 8'b11011011;
		20'b00010011000001110111: color_data = 8'b11011011;
		20'b00010011000001111000: color_data = 8'b11011011;
		20'b00010011000001111001: color_data = 8'b11011011;
		20'b00010011000001111010: color_data = 8'b11011011;
		20'b00010011000001111011: color_data = 8'b11011011;
		20'b00010011000001111100: color_data = 8'b11011011;
		20'b00010011000001111101: color_data = 8'b11011011;
		20'b00010011000001111110: color_data = 8'b11011011;
		20'b00010011000001111111: color_data = 8'b11011011;
		20'b00010011000010000000: color_data = 8'b11011011;
		20'b00010011000010000001: color_data = 8'b11011011;
		20'b00010011000010000010: color_data = 8'b11011011;
		20'b00010011000010000011: color_data = 8'b11011011;
		20'b00010011000010000100: color_data = 8'b11011011;
		20'b00010011000010000101: color_data = 8'b11011011;
		20'b00010011000010000110: color_data = 8'b11011011;
		20'b00010011000010000111: color_data = 8'b11011011;
		20'b00010011000010001000: color_data = 8'b11011011;
		20'b00010011000010001001: color_data = 8'b11011011;
		20'b00010011000010001010: color_data = 8'b11011011;
		20'b00010011000010001011: color_data = 8'b11011011;
		20'b00010011000010001100: color_data = 8'b11011011;
		20'b00010011000010001101: color_data = 8'b11011011;
		20'b00010011000010001110: color_data = 8'b11011011;
		20'b00010011000010011000: color_data = 8'b11011011;
		20'b00010011000010011001: color_data = 8'b11011011;
		20'b00010011000010011010: color_data = 8'b11011011;
		20'b00010011000010011011: color_data = 8'b11011011;
		20'b00010011000010011100: color_data = 8'b11011011;
		20'b00010011000010011101: color_data = 8'b11011011;
		20'b00010011000010011110: color_data = 8'b11011011;
		20'b00010011000010011111: color_data = 8'b11011011;
		20'b00010011000010100000: color_data = 8'b11011011;
		20'b00010011000010100001: color_data = 8'b11011011;
		20'b00010011000010100010: color_data = 8'b11011011;
		20'b00010011000010100011: color_data = 8'b11011011;
		20'b00010011000010100100: color_data = 8'b11011011;
		20'b00010011000010100101: color_data = 8'b11011011;
		20'b00010011000010100110: color_data = 8'b11011011;
		20'b00010011000010100111: color_data = 8'b11011011;
		20'b00010011000010101000: color_data = 8'b11011011;
		20'b00010011000010101001: color_data = 8'b11011011;
		20'b00010011000010101010: color_data = 8'b11011011;
		20'b00010011000010101011: color_data = 8'b11011011;
		20'b00010011000010101100: color_data = 8'b11011011;
		20'b00010011000010101101: color_data = 8'b11011011;
		20'b00010011000010101110: color_data = 8'b11011011;
		20'b00010011000010101111: color_data = 8'b11011011;
		20'b00010011000010110000: color_data = 8'b11011011;
		20'b00010011000010110001: color_data = 8'b11011011;
		20'b00010011000010110010: color_data = 8'b11011011;
		20'b00010011000010110011: color_data = 8'b11011011;
		20'b00010011000010110100: color_data = 8'b11011011;
		20'b00010011000010110101: color_data = 8'b11011011;
		20'b00010011000010110110: color_data = 8'b11011011;
		20'b00010011000010110111: color_data = 8'b11011011;
		20'b00010011000010111000: color_data = 8'b11011011;
		20'b00010011000010111001: color_data = 8'b11011011;
		20'b00010011000010111010: color_data = 8'b11011011;
		20'b00010011000010111011: color_data = 8'b11011011;
		20'b00010011000010111100: color_data = 8'b11011011;
		20'b00010011000010111101: color_data = 8'b11011011;
		20'b00010011000010111110: color_data = 8'b11011011;

		20'b00010011010000001001: color_data = 8'b11011011;
		20'b00010011010000001010: color_data = 8'b11111111;
		20'b00010011010000001011: color_data = 8'b11111111;
		20'b00010011010000001100: color_data = 8'b11111111;
		20'b00010011010000001101: color_data = 8'b11111111;
		20'b00010011010000001110: color_data = 8'b11111111;
		20'b00010011010000001111: color_data = 8'b11111111;
		20'b00010011010000010000: color_data = 8'b11111111;
		20'b00010011010000010001: color_data = 8'b11111111;
		20'b00010011010000010010: color_data = 8'b11111111;
		20'b00010011010000010011: color_data = 8'b11111111;
		20'b00010011010000010100: color_data = 8'b11111111;
		20'b00010011010000010101: color_data = 8'b11111111;
		20'b00010011010000010110: color_data = 8'b11111111;
		20'b00010011010000010111: color_data = 8'b11111111;
		20'b00010011010000011000: color_data = 8'b11111111;
		20'b00010011010000011001: color_data = 8'b11111111;
		20'b00010011010000011010: color_data = 8'b11111111;
		20'b00010011010000011011: color_data = 8'b11111111;
		20'b00010011010000011100: color_data = 8'b11111111;
		20'b00010011010000011101: color_data = 8'b11111111;
		20'b00010011010000011110: color_data = 8'b11111111;
		20'b00010011010000011111: color_data = 8'b11111111;
		20'b00010011010000100000: color_data = 8'b11111111;
		20'b00010011010000100001: color_data = 8'b11111111;
		20'b00010011010000100010: color_data = 8'b11111111;
		20'b00010011010000100011: color_data = 8'b11111111;
		20'b00010011010000100100: color_data = 8'b11111111;
		20'b00010011010000100101: color_data = 8'b11111111;
		20'b00010011010000100110: color_data = 8'b11111111;
		20'b00010011010000100111: color_data = 8'b11111111;
		20'b00010011010000101000: color_data = 8'b11111111;
		20'b00010011010000101001: color_data = 8'b11111111;
		20'b00010011010000101010: color_data = 8'b11111111;
		20'b00010011010000101011: color_data = 8'b11111111;
		20'b00010011010000101100: color_data = 8'b11111111;
		20'b00010011010000101101: color_data = 8'b11111111;
		20'b00010011010000101110: color_data = 8'b11111111;
		20'b00010011010000101111: color_data = 8'b11011011;
		20'b00010011010000111001: color_data = 8'b11111111;
		20'b00010011010000111010: color_data = 8'b11111111;
		20'b00010011010000111011: color_data = 8'b11111111;
		20'b00010011010000111100: color_data = 8'b11111111;
		20'b00010011010000111101: color_data = 8'b11111111;
		20'b00010011010000111110: color_data = 8'b11111111;
		20'b00010011010000111111: color_data = 8'b11111111;
		20'b00010011010001000000: color_data = 8'b11111111;
		20'b00010011010001000001: color_data = 8'b11111111;
		20'b00010011010001000010: color_data = 8'b11111111;
		20'b00010011010001000011: color_data = 8'b11111111;
		20'b00010011010001000100: color_data = 8'b11111111;
		20'b00010011010001000101: color_data = 8'b11111111;
		20'b00010011010001000110: color_data = 8'b11111111;
		20'b00010011010001000111: color_data = 8'b11111111;
		20'b00010011010001001000: color_data = 8'b11111111;
		20'b00010011010001001001: color_data = 8'b11111111;
		20'b00010011010001001010: color_data = 8'b11111111;
		20'b00010011010001001011: color_data = 8'b11111111;
		20'b00010011010001001100: color_data = 8'b11111111;
		20'b00010011010001001101: color_data = 8'b11111111;
		20'b00010011010001001110: color_data = 8'b11111111;
		20'b00010011010001001111: color_data = 8'b11111111;
		20'b00010011010001010000: color_data = 8'b11111111;
		20'b00010011010001010001: color_data = 8'b11111111;
		20'b00010011010001010010: color_data = 8'b11111111;
		20'b00010011010001010011: color_data = 8'b11111111;
		20'b00010011010001010100: color_data = 8'b11111111;
		20'b00010011010001010101: color_data = 8'b11111111;
		20'b00010011010001010110: color_data = 8'b11111111;
		20'b00010011010001010111: color_data = 8'b11111111;
		20'b00010011010001011000: color_data = 8'b11111111;
		20'b00010011010001011001: color_data = 8'b11111111;
		20'b00010011010001011010: color_data = 8'b11111111;
		20'b00010011010001011011: color_data = 8'b11111111;
		20'b00010011010001011100: color_data = 8'b11111111;
		20'b00010011010001011101: color_data = 8'b11111111;
		20'b00010011010001011110: color_data = 8'b11111111;
		20'b00010011010001011111: color_data = 8'b10010010;
		20'b00010011010001101000: color_data = 8'b10010010;
		20'b00010011010001101001: color_data = 8'b11111111;
		20'b00010011010001101010: color_data = 8'b11111111;
		20'b00010011010001101011: color_data = 8'b11111111;
		20'b00010011010001101100: color_data = 8'b11111111;
		20'b00010011010001101101: color_data = 8'b11111111;
		20'b00010011010001101110: color_data = 8'b11111111;
		20'b00010011010001101111: color_data = 8'b11111111;
		20'b00010011010001110000: color_data = 8'b11111111;
		20'b00010011010001110001: color_data = 8'b11111111;
		20'b00010011010001110010: color_data = 8'b11111111;
		20'b00010011010001110011: color_data = 8'b11111111;
		20'b00010011010001110100: color_data = 8'b11111111;
		20'b00010011010001110101: color_data = 8'b11111111;
		20'b00010011010001110110: color_data = 8'b11111111;
		20'b00010011010001110111: color_data = 8'b11111111;
		20'b00010011010001111000: color_data = 8'b11111111;
		20'b00010011010001111001: color_data = 8'b11111111;
		20'b00010011010001111010: color_data = 8'b11111111;
		20'b00010011010001111011: color_data = 8'b11111111;
		20'b00010011010001111100: color_data = 8'b11111111;
		20'b00010011010001111101: color_data = 8'b11111111;
		20'b00010011010001111110: color_data = 8'b11111111;
		20'b00010011010001111111: color_data = 8'b11111111;
		20'b00010011010010000000: color_data = 8'b11111111;
		20'b00010011010010000001: color_data = 8'b11111111;
		20'b00010011010010000010: color_data = 8'b11111111;
		20'b00010011010010000011: color_data = 8'b11111111;
		20'b00010011010010000100: color_data = 8'b11111111;
		20'b00010011010010000101: color_data = 8'b11111111;
		20'b00010011010010000110: color_data = 8'b11111111;
		20'b00010011010010000111: color_data = 8'b11111111;
		20'b00010011010010001000: color_data = 8'b11111111;
		20'b00010011010010001001: color_data = 8'b11111111;
		20'b00010011010010001010: color_data = 8'b11111111;
		20'b00010011010010001011: color_data = 8'b11111111;
		20'b00010011010010001100: color_data = 8'b11111111;
		20'b00010011010010001101: color_data = 8'b11111111;
		20'b00010011010010001110: color_data = 8'b11111111;
		20'b00010011010010011000: color_data = 8'b11011011;
		20'b00010011010010011001: color_data = 8'b11111111;
		20'b00010011010010011010: color_data = 8'b11111111;
		20'b00010011010010011011: color_data = 8'b11111111;
		20'b00010011010010011100: color_data = 8'b11111111;
		20'b00010011010010011101: color_data = 8'b11111111;
		20'b00010011010010011110: color_data = 8'b11111111;
		20'b00010011010010011111: color_data = 8'b11111111;
		20'b00010011010010100000: color_data = 8'b11111111;
		20'b00010011010010100001: color_data = 8'b11111111;
		20'b00010011010010100010: color_data = 8'b11111111;
		20'b00010011010010100011: color_data = 8'b11111111;
		20'b00010011010010100100: color_data = 8'b11111111;
		20'b00010011010010100101: color_data = 8'b11111111;
		20'b00010011010010100110: color_data = 8'b11111111;
		20'b00010011010010100111: color_data = 8'b11111111;
		20'b00010011010010101000: color_data = 8'b11111111;
		20'b00010011010010101001: color_data = 8'b11111111;
		20'b00010011010010101010: color_data = 8'b11111111;
		20'b00010011010010101011: color_data = 8'b11111111;
		20'b00010011010010101100: color_data = 8'b11111111;
		20'b00010011010010101101: color_data = 8'b11111111;
		20'b00010011010010101110: color_data = 8'b11111111;
		20'b00010011010010101111: color_data = 8'b11111111;
		20'b00010011010010110000: color_data = 8'b11111111;
		20'b00010011010010110001: color_data = 8'b11111111;
		20'b00010011010010110010: color_data = 8'b11111111;
		20'b00010011010010110011: color_data = 8'b11111111;
		20'b00010011010010110100: color_data = 8'b11111111;
		20'b00010011010010110101: color_data = 8'b11111111;
		20'b00010011010010110110: color_data = 8'b11111111;
		20'b00010011010010110111: color_data = 8'b11111111;
		20'b00010011010010111000: color_data = 8'b11111111;
		20'b00010011010010111001: color_data = 8'b11111111;
		20'b00010011010010111010: color_data = 8'b11111111;
		20'b00010011010010111011: color_data = 8'b11111111;
		20'b00010011010010111100: color_data = 8'b11111111;
		20'b00010011010010111101: color_data = 8'b11111111;
		20'b00010011010010111110: color_data = 8'b11011011;

		20'b00010011100000001001: color_data = 8'b11011011;
		20'b00010011100000001010: color_data = 8'b11111111;
		20'b00010011100000001011: color_data = 8'b11111111;
		20'b00010011100000001100: color_data = 8'b11111111;
		20'b00010011100000001101: color_data = 8'b11111111;
		20'b00010011100000001110: color_data = 8'b11111111;
		20'b00010011100000001111: color_data = 8'b11111111;
		20'b00010011100000010000: color_data = 8'b11111111;
		20'b00010011100000010001: color_data = 8'b11111111;
		20'b00010011100000010010: color_data = 8'b11111111;
		20'b00010011100000010011: color_data = 8'b11111111;
		20'b00010011100000010100: color_data = 8'b11111111;
		20'b00010011100000010101: color_data = 8'b11111111;
		20'b00010011100000010110: color_data = 8'b11111111;
		20'b00010011100000010111: color_data = 8'b11111111;
		20'b00010011100000011000: color_data = 8'b11111111;
		20'b00010011100000011001: color_data = 8'b11111111;
		20'b00010011100000011010: color_data = 8'b11111111;
		20'b00010011100000011011: color_data = 8'b11111111;
		20'b00010011100000011100: color_data = 8'b11111111;
		20'b00010011100000011101: color_data = 8'b11111111;
		20'b00010011100000011110: color_data = 8'b11111111;
		20'b00010011100000011111: color_data = 8'b11111111;
		20'b00010011100000100000: color_data = 8'b11111111;
		20'b00010011100000100001: color_data = 8'b11111111;
		20'b00010011100000100010: color_data = 8'b11111111;
		20'b00010011100000100011: color_data = 8'b11111111;
		20'b00010011100000100100: color_data = 8'b11111111;
		20'b00010011100000100101: color_data = 8'b11111111;
		20'b00010011100000100110: color_data = 8'b11111111;
		20'b00010011100000100111: color_data = 8'b11111111;
		20'b00010011100000101000: color_data = 8'b11111111;
		20'b00010011100000101001: color_data = 8'b11111111;
		20'b00010011100000101010: color_data = 8'b11111111;
		20'b00010011100000101011: color_data = 8'b11111111;
		20'b00010011100000101100: color_data = 8'b11111111;
		20'b00010011100000101101: color_data = 8'b11111111;
		20'b00010011100000101110: color_data = 8'b11111111;
		20'b00010011100000101111: color_data = 8'b11011011;
		20'b00010011100000111001: color_data = 8'b11111111;
		20'b00010011100000111010: color_data = 8'b11111111;
		20'b00010011100000111011: color_data = 8'b11111111;
		20'b00010011100000111100: color_data = 8'b11111111;
		20'b00010011100000111101: color_data = 8'b11111111;
		20'b00010011100000111110: color_data = 8'b11111111;
		20'b00010011100000111111: color_data = 8'b11111111;
		20'b00010011100001000000: color_data = 8'b11111111;
		20'b00010011100001000001: color_data = 8'b11111111;
		20'b00010011100001000010: color_data = 8'b11111111;
		20'b00010011100001000011: color_data = 8'b11111111;
		20'b00010011100001000100: color_data = 8'b11111111;
		20'b00010011100001000101: color_data = 8'b11111111;
		20'b00010011100001000110: color_data = 8'b11111111;
		20'b00010011100001000111: color_data = 8'b11111111;
		20'b00010011100001001000: color_data = 8'b11111111;
		20'b00010011100001001001: color_data = 8'b11111111;
		20'b00010011100001001010: color_data = 8'b11111111;
		20'b00010011100001001011: color_data = 8'b11111111;
		20'b00010011100001001100: color_data = 8'b11111111;
		20'b00010011100001001101: color_data = 8'b11111111;
		20'b00010011100001001110: color_data = 8'b11111111;
		20'b00010011100001001111: color_data = 8'b11111111;
		20'b00010011100001010000: color_data = 8'b11111111;
		20'b00010011100001010001: color_data = 8'b11111111;
		20'b00010011100001010010: color_data = 8'b11111111;
		20'b00010011100001010011: color_data = 8'b11111111;
		20'b00010011100001010100: color_data = 8'b11111111;
		20'b00010011100001010101: color_data = 8'b11111111;
		20'b00010011100001010110: color_data = 8'b11111111;
		20'b00010011100001010111: color_data = 8'b11111111;
		20'b00010011100001011000: color_data = 8'b11111111;
		20'b00010011100001011001: color_data = 8'b11111111;
		20'b00010011100001011010: color_data = 8'b11111111;
		20'b00010011100001011011: color_data = 8'b11111111;
		20'b00010011100001011100: color_data = 8'b11111111;
		20'b00010011100001011101: color_data = 8'b11111111;
		20'b00010011100001011110: color_data = 8'b11111111;
		20'b00010011100001011111: color_data = 8'b10010010;
		20'b00010011100001101000: color_data = 8'b10010010;
		20'b00010011100001101001: color_data = 8'b11111111;
		20'b00010011100001101010: color_data = 8'b11111111;
		20'b00010011100001101011: color_data = 8'b11111111;
		20'b00010011100001101100: color_data = 8'b11111111;
		20'b00010011100001101101: color_data = 8'b11111111;
		20'b00010011100001101110: color_data = 8'b11111111;
		20'b00010011100001101111: color_data = 8'b11111111;
		20'b00010011100001110000: color_data = 8'b11111111;
		20'b00010011100001110001: color_data = 8'b11111111;
		20'b00010011100001110010: color_data = 8'b11111111;
		20'b00010011100001110011: color_data = 8'b11111111;
		20'b00010011100001110100: color_data = 8'b11111111;
		20'b00010011100001110101: color_data = 8'b11111111;
		20'b00010011100001110110: color_data = 8'b11111111;
		20'b00010011100001110111: color_data = 8'b11111111;
		20'b00010011100001111000: color_data = 8'b11111111;
		20'b00010011100001111001: color_data = 8'b11111111;
		20'b00010011100001111010: color_data = 8'b11111111;
		20'b00010011100001111011: color_data = 8'b11111111;
		20'b00010011100001111100: color_data = 8'b11111111;
		20'b00010011100001111101: color_data = 8'b11111111;
		20'b00010011100001111110: color_data = 8'b11111111;
		20'b00010011100001111111: color_data = 8'b11111111;
		20'b00010011100010000000: color_data = 8'b11111111;
		20'b00010011100010000001: color_data = 8'b11111111;
		20'b00010011100010000010: color_data = 8'b11111111;
		20'b00010011100010000011: color_data = 8'b11111111;
		20'b00010011100010000100: color_data = 8'b11111111;
		20'b00010011100010000101: color_data = 8'b11111111;
		20'b00010011100010000110: color_data = 8'b11111111;
		20'b00010011100010000111: color_data = 8'b11111111;
		20'b00010011100010001000: color_data = 8'b11111111;
		20'b00010011100010001001: color_data = 8'b11111111;
		20'b00010011100010001010: color_data = 8'b11111111;
		20'b00010011100010001011: color_data = 8'b11111111;
		20'b00010011100010001100: color_data = 8'b11111111;
		20'b00010011100010001101: color_data = 8'b11111111;
		20'b00010011100010001110: color_data = 8'b11111111;
		20'b00010011100010011000: color_data = 8'b11011011;
		20'b00010011100010011001: color_data = 8'b11111111;
		20'b00010011100010011010: color_data = 8'b11111111;
		20'b00010011100010011011: color_data = 8'b11111111;
		20'b00010011100010011100: color_data = 8'b11111111;
		20'b00010011100010011101: color_data = 8'b11111111;
		20'b00010011100010011110: color_data = 8'b11111111;
		20'b00010011100010011111: color_data = 8'b11111111;
		20'b00010011100010100000: color_data = 8'b11111111;
		20'b00010011100010100001: color_data = 8'b11111111;
		20'b00010011100010100010: color_data = 8'b11111111;
		20'b00010011100010100011: color_data = 8'b11111111;
		20'b00010011100010100100: color_data = 8'b11111111;
		20'b00010011100010100101: color_data = 8'b11111111;
		20'b00010011100010100110: color_data = 8'b11111111;
		20'b00010011100010100111: color_data = 8'b11111111;
		20'b00010011100010101000: color_data = 8'b11111111;
		20'b00010011100010101001: color_data = 8'b11111111;
		20'b00010011100010101010: color_data = 8'b11111111;
		20'b00010011100010101011: color_data = 8'b11111111;
		20'b00010011100010101100: color_data = 8'b11111111;
		20'b00010011100010101101: color_data = 8'b11111111;
		20'b00010011100010101110: color_data = 8'b11111111;
		20'b00010011100010101111: color_data = 8'b11111111;
		20'b00010011100010110000: color_data = 8'b11111111;
		20'b00010011100010110001: color_data = 8'b11111111;
		20'b00010011100010110010: color_data = 8'b11111111;
		20'b00010011100010110011: color_data = 8'b11111111;
		20'b00010011100010110100: color_data = 8'b11111111;
		20'b00010011100010110101: color_data = 8'b11111111;
		20'b00010011100010110110: color_data = 8'b11111111;
		20'b00010011100010110111: color_data = 8'b11111111;
		20'b00010011100010111000: color_data = 8'b11111111;
		20'b00010011100010111001: color_data = 8'b11111111;
		20'b00010011100010111010: color_data = 8'b11111111;
		20'b00010011100010111011: color_data = 8'b11111111;
		20'b00010011100010111100: color_data = 8'b11111111;
		20'b00010011100010111101: color_data = 8'b11111111;
		20'b00010011100010111110: color_data = 8'b11011011;

		20'b00010011110000001001: color_data = 8'b11011011;
		20'b00010011110000001010: color_data = 8'b11111111;
		20'b00010011110000001011: color_data = 8'b11111111;
		20'b00010011110000001100: color_data = 8'b11111111;
		20'b00010011110000001101: color_data = 8'b11111111;
		20'b00010011110000001110: color_data = 8'b11111111;
		20'b00010011110000001111: color_data = 8'b11111111;
		20'b00010011110000010000: color_data = 8'b11111111;
		20'b00010011110000010001: color_data = 8'b11111111;
		20'b00010011110000010010: color_data = 8'b11111111;
		20'b00010011110000010011: color_data = 8'b11111111;
		20'b00010011110000010100: color_data = 8'b11111111;
		20'b00010011110000010101: color_data = 8'b11111111;
		20'b00010011110000010110: color_data = 8'b11111111;
		20'b00010011110000010111: color_data = 8'b11111111;
		20'b00010011110000011000: color_data = 8'b11111111;
		20'b00010011110000011001: color_data = 8'b11111111;
		20'b00010011110000011010: color_data = 8'b11111111;
		20'b00010011110000011011: color_data = 8'b11111111;
		20'b00010011110000011100: color_data = 8'b11111111;
		20'b00010011110000011101: color_data = 8'b11111111;
		20'b00010011110000011110: color_data = 8'b11111111;
		20'b00010011110000011111: color_data = 8'b11111111;
		20'b00010011110000100000: color_data = 8'b11111111;
		20'b00010011110000100001: color_data = 8'b11111111;
		20'b00010011110000100010: color_data = 8'b11111111;
		20'b00010011110000100011: color_data = 8'b11111111;
		20'b00010011110000100100: color_data = 8'b11111111;
		20'b00010011110000100101: color_data = 8'b11111111;
		20'b00010011110000100110: color_data = 8'b11111111;
		20'b00010011110000100111: color_data = 8'b11111111;
		20'b00010011110000101000: color_data = 8'b11111111;
		20'b00010011110000101001: color_data = 8'b11111111;
		20'b00010011110000101010: color_data = 8'b11111111;
		20'b00010011110000101011: color_data = 8'b11111111;
		20'b00010011110000101100: color_data = 8'b11111111;
		20'b00010011110000101101: color_data = 8'b11111111;
		20'b00010011110000101110: color_data = 8'b11111111;
		20'b00010011110000101111: color_data = 8'b11011011;
		20'b00010011110000111001: color_data = 8'b11111111;
		20'b00010011110000111010: color_data = 8'b11111111;
		20'b00010011110000111011: color_data = 8'b11111111;
		20'b00010011110000111100: color_data = 8'b11111111;
		20'b00010011110000111101: color_data = 8'b11111111;
		20'b00010011110000111110: color_data = 8'b11111111;
		20'b00010011110000111111: color_data = 8'b11111111;
		20'b00010011110001000000: color_data = 8'b11111111;
		20'b00010011110001000001: color_data = 8'b11111111;
		20'b00010011110001000010: color_data = 8'b11111111;
		20'b00010011110001000011: color_data = 8'b11111111;
		20'b00010011110001000100: color_data = 8'b11111111;
		20'b00010011110001000101: color_data = 8'b11111111;
		20'b00010011110001000110: color_data = 8'b11111111;
		20'b00010011110001000111: color_data = 8'b11111111;
		20'b00010011110001001000: color_data = 8'b11111111;
		20'b00010011110001001001: color_data = 8'b11111111;
		20'b00010011110001001010: color_data = 8'b11111111;
		20'b00010011110001001011: color_data = 8'b11111111;
		20'b00010011110001001100: color_data = 8'b11111111;
		20'b00010011110001001101: color_data = 8'b11111111;
		20'b00010011110001001110: color_data = 8'b11111111;
		20'b00010011110001001111: color_data = 8'b11111111;
		20'b00010011110001010000: color_data = 8'b11111111;
		20'b00010011110001010001: color_data = 8'b11111111;
		20'b00010011110001010010: color_data = 8'b11111111;
		20'b00010011110001010011: color_data = 8'b11111111;
		20'b00010011110001010100: color_data = 8'b11111111;
		20'b00010011110001010101: color_data = 8'b11111111;
		20'b00010011110001010110: color_data = 8'b11111111;
		20'b00010011110001010111: color_data = 8'b11111111;
		20'b00010011110001011000: color_data = 8'b11111111;
		20'b00010011110001011001: color_data = 8'b11111111;
		20'b00010011110001011010: color_data = 8'b11111111;
		20'b00010011110001011011: color_data = 8'b11111111;
		20'b00010011110001011100: color_data = 8'b11111111;
		20'b00010011110001011101: color_data = 8'b11111111;
		20'b00010011110001011110: color_data = 8'b11111111;
		20'b00010011110001011111: color_data = 8'b10010010;
		20'b00010011110001101000: color_data = 8'b10010010;
		20'b00010011110001101001: color_data = 8'b11111111;
		20'b00010011110001101010: color_data = 8'b11111111;
		20'b00010011110001101011: color_data = 8'b11111111;
		20'b00010011110001101100: color_data = 8'b11111111;
		20'b00010011110001101101: color_data = 8'b11111111;
		20'b00010011110001101110: color_data = 8'b11111111;
		20'b00010011110001101111: color_data = 8'b11111111;
		20'b00010011110001110000: color_data = 8'b11111111;
		20'b00010011110001110001: color_data = 8'b11111111;
		20'b00010011110001110010: color_data = 8'b11111111;
		20'b00010011110001110011: color_data = 8'b11111111;
		20'b00010011110001110100: color_data = 8'b11111111;
		20'b00010011110001110101: color_data = 8'b11111111;
		20'b00010011110001110110: color_data = 8'b11111111;
		20'b00010011110001110111: color_data = 8'b11111111;
		20'b00010011110001111000: color_data = 8'b11111111;
		20'b00010011110001111001: color_data = 8'b11111111;
		20'b00010011110001111010: color_data = 8'b11111111;
		20'b00010011110001111011: color_data = 8'b11111111;
		20'b00010011110001111100: color_data = 8'b11111111;
		20'b00010011110001111101: color_data = 8'b11111111;
		20'b00010011110001111110: color_data = 8'b11111111;
		20'b00010011110001111111: color_data = 8'b11111111;
		20'b00010011110010000000: color_data = 8'b11111111;
		20'b00010011110010000001: color_data = 8'b11111111;
		20'b00010011110010000010: color_data = 8'b11111111;
		20'b00010011110010000011: color_data = 8'b11111111;
		20'b00010011110010000100: color_data = 8'b11111111;
		20'b00010011110010000101: color_data = 8'b11111111;
		20'b00010011110010000110: color_data = 8'b11111111;
		20'b00010011110010000111: color_data = 8'b11111111;
		20'b00010011110010001000: color_data = 8'b11111111;
		20'b00010011110010001001: color_data = 8'b11111111;
		20'b00010011110010001010: color_data = 8'b11111111;
		20'b00010011110010001011: color_data = 8'b11111111;
		20'b00010011110010001100: color_data = 8'b11111111;
		20'b00010011110010001101: color_data = 8'b11111111;
		20'b00010011110010001110: color_data = 8'b11111111;
		20'b00010011110010011000: color_data = 8'b11011011;
		20'b00010011110010011001: color_data = 8'b11111111;
		20'b00010011110010011010: color_data = 8'b11111111;
		20'b00010011110010011011: color_data = 8'b11111111;
		20'b00010011110010011100: color_data = 8'b11111111;
		20'b00010011110010011101: color_data = 8'b11111111;
		20'b00010011110010011110: color_data = 8'b11111111;
		20'b00010011110010011111: color_data = 8'b11111111;
		20'b00010011110010100000: color_data = 8'b11111111;
		20'b00010011110010100001: color_data = 8'b11111111;
		20'b00010011110010100010: color_data = 8'b11111111;
		20'b00010011110010100011: color_data = 8'b11111111;
		20'b00010011110010100100: color_data = 8'b11111111;
		20'b00010011110010100101: color_data = 8'b11111111;
		20'b00010011110010100110: color_data = 8'b11111111;
		20'b00010011110010100111: color_data = 8'b11111111;
		20'b00010011110010101000: color_data = 8'b11111111;
		20'b00010011110010101001: color_data = 8'b11111111;
		20'b00010011110010101010: color_data = 8'b11111111;
		20'b00010011110010101011: color_data = 8'b11111111;
		20'b00010011110010101100: color_data = 8'b11111111;
		20'b00010011110010101101: color_data = 8'b11111111;
		20'b00010011110010101110: color_data = 8'b11111111;
		20'b00010011110010101111: color_data = 8'b11111111;
		20'b00010011110010110000: color_data = 8'b11111111;
		20'b00010011110010110001: color_data = 8'b11111111;
		20'b00010011110010110010: color_data = 8'b11111111;
		20'b00010011110010110011: color_data = 8'b11111111;
		20'b00010011110010110100: color_data = 8'b11111111;
		20'b00010011110010110101: color_data = 8'b11111111;
		20'b00010011110010110110: color_data = 8'b11111111;
		20'b00010011110010110111: color_data = 8'b11111111;
		20'b00010011110010111000: color_data = 8'b11111111;
		20'b00010011110010111001: color_data = 8'b11111111;
		20'b00010011110010111010: color_data = 8'b11111111;
		20'b00010011110010111011: color_data = 8'b11111111;
		20'b00010011110010111100: color_data = 8'b11111111;
		20'b00010011110010111101: color_data = 8'b11111111;
		20'b00010011110010111110: color_data = 8'b11011011;

		20'b00010100000000001001: color_data = 8'b11011011;
		20'b00010100000000001010: color_data = 8'b11111111;
		20'b00010100000000001011: color_data = 8'b11111111;
		20'b00010100000000001100: color_data = 8'b11111111;
		20'b00010100000000001101: color_data = 8'b11111111;
		20'b00010100000000001110: color_data = 8'b11111111;
		20'b00010100000000001111: color_data = 8'b11111111;
		20'b00010100000000010000: color_data = 8'b11111111;
		20'b00010100000000010001: color_data = 8'b11111111;
		20'b00010100000000010010: color_data = 8'b11111111;
		20'b00010100000000010011: color_data = 8'b11111111;
		20'b00010100000000010100: color_data = 8'b11111111;
		20'b00010100000000010101: color_data = 8'b11111111;
		20'b00010100000000010110: color_data = 8'b11111111;
		20'b00010100000000010111: color_data = 8'b11111111;
		20'b00010100000000011000: color_data = 8'b11111111;
		20'b00010100000000011001: color_data = 8'b11111111;
		20'b00010100000000011010: color_data = 8'b11111111;
		20'b00010100000000011011: color_data = 8'b11111111;
		20'b00010100000000011100: color_data = 8'b11111111;
		20'b00010100000000011101: color_data = 8'b11111111;
		20'b00010100000000011110: color_data = 8'b11111111;
		20'b00010100000000011111: color_data = 8'b11111111;
		20'b00010100000000100000: color_data = 8'b11111111;
		20'b00010100000000100001: color_data = 8'b11111111;
		20'b00010100000000100010: color_data = 8'b11111111;
		20'b00010100000000100011: color_data = 8'b11111111;
		20'b00010100000000100100: color_data = 8'b11111111;
		20'b00010100000000100101: color_data = 8'b11111111;
		20'b00010100000000100110: color_data = 8'b11111111;
		20'b00010100000000100111: color_data = 8'b11111111;
		20'b00010100000000101000: color_data = 8'b11111111;
		20'b00010100000000101001: color_data = 8'b11111111;
		20'b00010100000000101010: color_data = 8'b11111111;
		20'b00010100000000101011: color_data = 8'b11111111;
		20'b00010100000000101100: color_data = 8'b11111111;
		20'b00010100000000101101: color_data = 8'b11111111;
		20'b00010100000000101110: color_data = 8'b11111111;
		20'b00010100000000101111: color_data = 8'b11011011;
		20'b00010100000000111001: color_data = 8'b11111111;
		20'b00010100000000111010: color_data = 8'b11111111;
		20'b00010100000000111011: color_data = 8'b11111111;
		20'b00010100000000111100: color_data = 8'b11111111;
		20'b00010100000000111101: color_data = 8'b11111111;
		20'b00010100000000111110: color_data = 8'b11111111;
		20'b00010100000000111111: color_data = 8'b11111111;
		20'b00010100000001000000: color_data = 8'b11111111;
		20'b00010100000001000001: color_data = 8'b11111111;
		20'b00010100000001000010: color_data = 8'b11111111;
		20'b00010100000001000011: color_data = 8'b11111111;
		20'b00010100000001000100: color_data = 8'b11111111;
		20'b00010100000001000101: color_data = 8'b11111111;
		20'b00010100000001000110: color_data = 8'b11111111;
		20'b00010100000001000111: color_data = 8'b11111111;
		20'b00010100000001001000: color_data = 8'b11111111;
		20'b00010100000001001001: color_data = 8'b11111111;
		20'b00010100000001001010: color_data = 8'b11111111;
		20'b00010100000001001011: color_data = 8'b11111111;
		20'b00010100000001001100: color_data = 8'b11111111;
		20'b00010100000001001101: color_data = 8'b11111111;
		20'b00010100000001001110: color_data = 8'b11111111;
		20'b00010100000001001111: color_data = 8'b11111111;
		20'b00010100000001010000: color_data = 8'b11111111;
		20'b00010100000001010001: color_data = 8'b11111111;
		20'b00010100000001010010: color_data = 8'b11111111;
		20'b00010100000001010011: color_data = 8'b11111111;
		20'b00010100000001010100: color_data = 8'b11111111;
		20'b00010100000001010101: color_data = 8'b11111111;
		20'b00010100000001010110: color_data = 8'b11111111;
		20'b00010100000001010111: color_data = 8'b11111111;
		20'b00010100000001011000: color_data = 8'b11111111;
		20'b00010100000001011001: color_data = 8'b11111111;
		20'b00010100000001011010: color_data = 8'b11111111;
		20'b00010100000001011011: color_data = 8'b11111111;
		20'b00010100000001011100: color_data = 8'b11111111;
		20'b00010100000001011101: color_data = 8'b11111111;
		20'b00010100000001011110: color_data = 8'b11111111;
		20'b00010100000001011111: color_data = 8'b10010010;
		20'b00010100000001101000: color_data = 8'b10010010;
		20'b00010100000001101001: color_data = 8'b11111111;
		20'b00010100000001101010: color_data = 8'b11111111;
		20'b00010100000001101011: color_data = 8'b11111111;
		20'b00010100000001101100: color_data = 8'b11111111;
		20'b00010100000001101101: color_data = 8'b11111111;
		20'b00010100000001101110: color_data = 8'b11111111;
		20'b00010100000001101111: color_data = 8'b11111111;
		20'b00010100000001110000: color_data = 8'b11111111;
		20'b00010100000001110001: color_data = 8'b11111111;
		20'b00010100000001110010: color_data = 8'b11111111;
		20'b00010100000001110011: color_data = 8'b11111111;
		20'b00010100000001110100: color_data = 8'b11111111;
		20'b00010100000001110101: color_data = 8'b11111111;
		20'b00010100000001110110: color_data = 8'b11111111;
		20'b00010100000001110111: color_data = 8'b11111111;
		20'b00010100000001111000: color_data = 8'b11111111;
		20'b00010100000001111001: color_data = 8'b11111111;
		20'b00010100000001111010: color_data = 8'b11111111;
		20'b00010100000001111011: color_data = 8'b11111111;
		20'b00010100000001111100: color_data = 8'b11111111;
		20'b00010100000001111101: color_data = 8'b11111111;
		20'b00010100000001111110: color_data = 8'b11111111;
		20'b00010100000001111111: color_data = 8'b11111111;
		20'b00010100000010000000: color_data = 8'b11111111;
		20'b00010100000010000001: color_data = 8'b11111111;
		20'b00010100000010000010: color_data = 8'b11111111;
		20'b00010100000010000011: color_data = 8'b11111111;
		20'b00010100000010000100: color_data = 8'b11111111;
		20'b00010100000010000101: color_data = 8'b11111111;
		20'b00010100000010000110: color_data = 8'b11111111;
		20'b00010100000010000111: color_data = 8'b11111111;
		20'b00010100000010001000: color_data = 8'b11111111;
		20'b00010100000010001001: color_data = 8'b11111111;
		20'b00010100000010001010: color_data = 8'b11111111;
		20'b00010100000010001011: color_data = 8'b11111111;
		20'b00010100000010001100: color_data = 8'b11111111;
		20'b00010100000010001101: color_data = 8'b11111111;
		20'b00010100000010001110: color_data = 8'b11111111;
		20'b00010100000010011000: color_data = 8'b11011011;
		20'b00010100000010011001: color_data = 8'b11111111;
		20'b00010100000010011010: color_data = 8'b11111111;
		20'b00010100000010011011: color_data = 8'b11111111;
		20'b00010100000010011100: color_data = 8'b11111111;
		20'b00010100000010011101: color_data = 8'b11111111;
		20'b00010100000010011110: color_data = 8'b11111111;
		20'b00010100000010011111: color_data = 8'b11111111;
		20'b00010100000010100000: color_data = 8'b11111111;
		20'b00010100000010100001: color_data = 8'b11111111;
		20'b00010100000010100010: color_data = 8'b11111111;
		20'b00010100000010100011: color_data = 8'b11111111;
		20'b00010100000010100100: color_data = 8'b11111111;
		20'b00010100000010100101: color_data = 8'b11111111;
		20'b00010100000010100110: color_data = 8'b11111111;
		20'b00010100000010100111: color_data = 8'b11111111;
		20'b00010100000010101000: color_data = 8'b11111111;
		20'b00010100000010101001: color_data = 8'b11111111;
		20'b00010100000010101010: color_data = 8'b11111111;
		20'b00010100000010101011: color_data = 8'b11111111;
		20'b00010100000010101100: color_data = 8'b11111111;
		20'b00010100000010101101: color_data = 8'b11111111;
		20'b00010100000010101110: color_data = 8'b11111111;
		20'b00010100000010101111: color_data = 8'b11111111;
		20'b00010100000010110000: color_data = 8'b11111111;
		20'b00010100000010110001: color_data = 8'b11111111;
		20'b00010100000010110010: color_data = 8'b11111111;
		20'b00010100000010110011: color_data = 8'b11111111;
		20'b00010100000010110100: color_data = 8'b11111111;
		20'b00010100000010110101: color_data = 8'b11111111;
		20'b00010100000010110110: color_data = 8'b11111111;
		20'b00010100000010110111: color_data = 8'b11111111;
		20'b00010100000010111000: color_data = 8'b11111111;
		20'b00010100000010111001: color_data = 8'b11111111;
		20'b00010100000010111010: color_data = 8'b11111111;
		20'b00010100000010111011: color_data = 8'b11111111;
		20'b00010100000010111100: color_data = 8'b11111111;
		20'b00010100000010111101: color_data = 8'b11111111;
		20'b00010100000010111110: color_data = 8'b11011011;

		20'b00010100010000001001: color_data = 8'b11011011;
		20'b00010100010000001010: color_data = 8'b11111111;
		20'b00010100010000001011: color_data = 8'b11111111;
		20'b00010100010000001100: color_data = 8'b11111111;
		20'b00010100010000001101: color_data = 8'b11111111;
		20'b00010100010000001110: color_data = 8'b11111111;
		20'b00010100010000001111: color_data = 8'b11111111;
		20'b00010100010000010000: color_data = 8'b11111111;
		20'b00010100010000010001: color_data = 8'b11111111;
		20'b00010100010000010010: color_data = 8'b11111111;
		20'b00010100010000010011: color_data = 8'b11111111;
		20'b00010100010000010100: color_data = 8'b11111111;
		20'b00010100010000010101: color_data = 8'b11111111;
		20'b00010100010000010110: color_data = 8'b11111111;
		20'b00010100010000010111: color_data = 8'b11111111;
		20'b00010100010000011000: color_data = 8'b11111111;
		20'b00010100010000011001: color_data = 8'b11111111;
		20'b00010100010000011010: color_data = 8'b11111111;
		20'b00010100010000011011: color_data = 8'b11111111;
		20'b00010100010000011100: color_data = 8'b11111111;
		20'b00010100010000011101: color_data = 8'b11111111;
		20'b00010100010000011110: color_data = 8'b11111111;
		20'b00010100010000011111: color_data = 8'b11111111;
		20'b00010100010000100000: color_data = 8'b11111111;
		20'b00010100010000100001: color_data = 8'b11111111;
		20'b00010100010000100010: color_data = 8'b11111111;
		20'b00010100010000100011: color_data = 8'b11111111;
		20'b00010100010000100100: color_data = 8'b11111111;
		20'b00010100010000100101: color_data = 8'b11111111;
		20'b00010100010000100110: color_data = 8'b11111111;
		20'b00010100010000100111: color_data = 8'b11111111;
		20'b00010100010000101000: color_data = 8'b11111111;
		20'b00010100010000101001: color_data = 8'b11111111;
		20'b00010100010000101010: color_data = 8'b11111111;
		20'b00010100010000101011: color_data = 8'b11111111;
		20'b00010100010000101100: color_data = 8'b11111111;
		20'b00010100010000101101: color_data = 8'b11111111;
		20'b00010100010000101110: color_data = 8'b11111111;
		20'b00010100010000101111: color_data = 8'b11011011;
		20'b00010100010000111001: color_data = 8'b11111111;
		20'b00010100010000111010: color_data = 8'b11111111;
		20'b00010100010000111011: color_data = 8'b11111111;
		20'b00010100010000111100: color_data = 8'b11111111;
		20'b00010100010000111101: color_data = 8'b11111111;
		20'b00010100010000111110: color_data = 8'b11111111;
		20'b00010100010000111111: color_data = 8'b11111111;
		20'b00010100010001000000: color_data = 8'b11111111;
		20'b00010100010001000001: color_data = 8'b11111111;
		20'b00010100010001000010: color_data = 8'b11111111;
		20'b00010100010001000011: color_data = 8'b11111111;
		20'b00010100010001000100: color_data = 8'b11111111;
		20'b00010100010001000101: color_data = 8'b11111111;
		20'b00010100010001000110: color_data = 8'b11111111;
		20'b00010100010001000111: color_data = 8'b11111111;
		20'b00010100010001001000: color_data = 8'b11111111;
		20'b00010100010001001001: color_data = 8'b11111111;
		20'b00010100010001001010: color_data = 8'b11111111;
		20'b00010100010001001011: color_data = 8'b11111111;
		20'b00010100010001001100: color_data = 8'b11111111;
		20'b00010100010001001101: color_data = 8'b11111111;
		20'b00010100010001001110: color_data = 8'b11111111;
		20'b00010100010001001111: color_data = 8'b11111111;
		20'b00010100010001010000: color_data = 8'b11111111;
		20'b00010100010001010001: color_data = 8'b11111111;
		20'b00010100010001010010: color_data = 8'b11111111;
		20'b00010100010001010011: color_data = 8'b11111111;
		20'b00010100010001010100: color_data = 8'b11111111;
		20'b00010100010001010101: color_data = 8'b11111111;
		20'b00010100010001010110: color_data = 8'b11111111;
		20'b00010100010001010111: color_data = 8'b11111111;
		20'b00010100010001011000: color_data = 8'b11111111;
		20'b00010100010001011001: color_data = 8'b11111111;
		20'b00010100010001011010: color_data = 8'b11111111;
		20'b00010100010001011011: color_data = 8'b11111111;
		20'b00010100010001011100: color_data = 8'b11111111;
		20'b00010100010001011101: color_data = 8'b11111111;
		20'b00010100010001011110: color_data = 8'b11111111;
		20'b00010100010001011111: color_data = 8'b10010010;
		20'b00010100010001101000: color_data = 8'b10010010;
		20'b00010100010001101001: color_data = 8'b11111111;
		20'b00010100010001101010: color_data = 8'b11111111;
		20'b00010100010001101011: color_data = 8'b11111111;
		20'b00010100010001101100: color_data = 8'b11111111;
		20'b00010100010001101101: color_data = 8'b11111111;
		20'b00010100010001101110: color_data = 8'b11111111;
		20'b00010100010001101111: color_data = 8'b11111111;
		20'b00010100010001110000: color_data = 8'b11111111;
		20'b00010100010001110001: color_data = 8'b11111111;
		20'b00010100010001110010: color_data = 8'b11111111;
		20'b00010100010001110011: color_data = 8'b11111111;
		20'b00010100010001110100: color_data = 8'b11111111;
		20'b00010100010001110101: color_data = 8'b11111111;
		20'b00010100010001110110: color_data = 8'b11111111;
		20'b00010100010001110111: color_data = 8'b11111111;
		20'b00010100010001111000: color_data = 8'b11111111;
		20'b00010100010001111001: color_data = 8'b11111111;
		20'b00010100010001111010: color_data = 8'b11111111;
		20'b00010100010001111011: color_data = 8'b11111111;
		20'b00010100010001111100: color_data = 8'b11111111;
		20'b00010100010001111101: color_data = 8'b11111111;
		20'b00010100010001111110: color_data = 8'b11111111;
		20'b00010100010001111111: color_data = 8'b11111111;
		20'b00010100010010000000: color_data = 8'b11111111;
		20'b00010100010010000001: color_data = 8'b11111111;
		20'b00010100010010000010: color_data = 8'b11111111;
		20'b00010100010010000011: color_data = 8'b11111111;
		20'b00010100010010000100: color_data = 8'b11111111;
		20'b00010100010010000101: color_data = 8'b11111111;
		20'b00010100010010000110: color_data = 8'b11111111;
		20'b00010100010010000111: color_data = 8'b11111111;
		20'b00010100010010001000: color_data = 8'b11111111;
		20'b00010100010010001001: color_data = 8'b11111111;
		20'b00010100010010001010: color_data = 8'b11111111;
		20'b00010100010010001011: color_data = 8'b11111111;
		20'b00010100010010001100: color_data = 8'b11111111;
		20'b00010100010010001101: color_data = 8'b11111111;
		20'b00010100010010001110: color_data = 8'b11111111;
		20'b00010100010010011000: color_data = 8'b11011011;
		20'b00010100010010011001: color_data = 8'b11111111;
		20'b00010100010010011010: color_data = 8'b11111111;
		20'b00010100010010011011: color_data = 8'b11111111;
		20'b00010100010010011100: color_data = 8'b11111111;
		20'b00010100010010011101: color_data = 8'b11111111;
		20'b00010100010010011110: color_data = 8'b11111111;
		20'b00010100010010011111: color_data = 8'b11111111;
		20'b00010100010010100000: color_data = 8'b11111111;
		20'b00010100010010100001: color_data = 8'b11111111;
		20'b00010100010010100010: color_data = 8'b11111111;
		20'b00010100010010100011: color_data = 8'b11111111;
		20'b00010100010010100100: color_data = 8'b11111111;
		20'b00010100010010100101: color_data = 8'b11111111;
		20'b00010100010010100110: color_data = 8'b11111111;
		20'b00010100010010100111: color_data = 8'b11111111;
		20'b00010100010010101000: color_data = 8'b11111111;
		20'b00010100010010101001: color_data = 8'b11111111;
		20'b00010100010010101010: color_data = 8'b11111111;
		20'b00010100010010101011: color_data = 8'b11111111;
		20'b00010100010010101100: color_data = 8'b11111111;
		20'b00010100010010101101: color_data = 8'b11111111;
		20'b00010100010010101110: color_data = 8'b11111111;
		20'b00010100010010101111: color_data = 8'b11111111;
		20'b00010100010010110000: color_data = 8'b11111111;
		20'b00010100010010110001: color_data = 8'b11111111;
		20'b00010100010010110010: color_data = 8'b11111111;
		20'b00010100010010110011: color_data = 8'b11111111;
		20'b00010100010010110100: color_data = 8'b11111111;
		20'b00010100010010110101: color_data = 8'b11111111;
		20'b00010100010010110110: color_data = 8'b11111111;
		20'b00010100010010110111: color_data = 8'b11111111;
		20'b00010100010010111000: color_data = 8'b11111111;
		20'b00010100010010111001: color_data = 8'b11111111;
		20'b00010100010010111010: color_data = 8'b11111111;
		20'b00010100010010111011: color_data = 8'b11111111;
		20'b00010100010010111100: color_data = 8'b11111111;
		20'b00010100010010111101: color_data = 8'b11111111;
		20'b00010100010010111110: color_data = 8'b11011011;

		20'b00010100100000001001: color_data = 8'b11011011;
		20'b00010100100000001010: color_data = 8'b11111111;
		20'b00010100100000001011: color_data = 8'b11111111;
		20'b00010100100000001100: color_data = 8'b11111111;
		20'b00010100100000001101: color_data = 8'b11111111;
		20'b00010100100000001110: color_data = 8'b11111111;
		20'b00010100100000001111: color_data = 8'b11111111;
		20'b00010100100000010000: color_data = 8'b11111111;
		20'b00010100100000010001: color_data = 8'b11111111;
		20'b00010100100000010010: color_data = 8'b11111111;
		20'b00010100100000010011: color_data = 8'b11111111;
		20'b00010100100000010100: color_data = 8'b11111111;
		20'b00010100100000010101: color_data = 8'b11111111;
		20'b00010100100000010110: color_data = 8'b11111111;
		20'b00010100100000010111: color_data = 8'b11111111;
		20'b00010100100000011000: color_data = 8'b11111111;
		20'b00010100100000011001: color_data = 8'b11111111;
		20'b00010100100000011010: color_data = 8'b11111111;
		20'b00010100100000011011: color_data = 8'b11111111;
		20'b00010100100000011100: color_data = 8'b11111111;
		20'b00010100100000011101: color_data = 8'b11111111;
		20'b00010100100000011110: color_data = 8'b11111111;
		20'b00010100100000011111: color_data = 8'b11111111;
		20'b00010100100000100000: color_data = 8'b11111111;
		20'b00010100100000100001: color_data = 8'b11111111;
		20'b00010100100000100010: color_data = 8'b11111111;
		20'b00010100100000100011: color_data = 8'b11111111;
		20'b00010100100000100100: color_data = 8'b11111111;
		20'b00010100100000100101: color_data = 8'b11111111;
		20'b00010100100000100110: color_data = 8'b11111111;
		20'b00010100100000100111: color_data = 8'b11111111;
		20'b00010100100000101000: color_data = 8'b11111111;
		20'b00010100100000101001: color_data = 8'b11111111;
		20'b00010100100000101010: color_data = 8'b11111111;
		20'b00010100100000101011: color_data = 8'b11111111;
		20'b00010100100000101100: color_data = 8'b11111111;
		20'b00010100100000101101: color_data = 8'b11111111;
		20'b00010100100000101110: color_data = 8'b11111111;
		20'b00010100100000101111: color_data = 8'b11011011;
		20'b00010100100000111001: color_data = 8'b11111111;
		20'b00010100100000111010: color_data = 8'b11111111;
		20'b00010100100000111011: color_data = 8'b11111111;
		20'b00010100100000111100: color_data = 8'b11111111;
		20'b00010100100000111101: color_data = 8'b11111111;
		20'b00010100100000111110: color_data = 8'b11111111;
		20'b00010100100000111111: color_data = 8'b11111111;
		20'b00010100100001000000: color_data = 8'b11111111;
		20'b00010100100001000001: color_data = 8'b11111111;
		20'b00010100100001000010: color_data = 8'b11111111;
		20'b00010100100001000011: color_data = 8'b11111111;
		20'b00010100100001000100: color_data = 8'b11111111;
		20'b00010100100001000101: color_data = 8'b11111111;
		20'b00010100100001000110: color_data = 8'b11111111;
		20'b00010100100001000111: color_data = 8'b11111111;
		20'b00010100100001001000: color_data = 8'b11111111;
		20'b00010100100001001001: color_data = 8'b11111111;
		20'b00010100100001001010: color_data = 8'b11111111;
		20'b00010100100001001011: color_data = 8'b11111111;
		20'b00010100100001001100: color_data = 8'b11111111;
		20'b00010100100001001101: color_data = 8'b11111111;
		20'b00010100100001001110: color_data = 8'b11111111;
		20'b00010100100001001111: color_data = 8'b11111111;
		20'b00010100100001010000: color_data = 8'b11111111;
		20'b00010100100001010001: color_data = 8'b11111111;
		20'b00010100100001010010: color_data = 8'b11111111;
		20'b00010100100001010011: color_data = 8'b11111111;
		20'b00010100100001010100: color_data = 8'b11111111;
		20'b00010100100001010101: color_data = 8'b11111111;
		20'b00010100100001010110: color_data = 8'b11111111;
		20'b00010100100001010111: color_data = 8'b11111111;
		20'b00010100100001011000: color_data = 8'b11111111;
		20'b00010100100001011001: color_data = 8'b11111111;
		20'b00010100100001011010: color_data = 8'b11111111;
		20'b00010100100001011011: color_data = 8'b11111111;
		20'b00010100100001011100: color_data = 8'b11111111;
		20'b00010100100001011101: color_data = 8'b11111111;
		20'b00010100100001011110: color_data = 8'b11111111;
		20'b00010100100001011111: color_data = 8'b10010010;
		20'b00010100100001101000: color_data = 8'b10010010;
		20'b00010100100001101001: color_data = 8'b11111111;
		20'b00010100100001101010: color_data = 8'b11111111;
		20'b00010100100001101011: color_data = 8'b11111111;
		20'b00010100100001101100: color_data = 8'b11111111;
		20'b00010100100001101101: color_data = 8'b11111111;
		20'b00010100100001101110: color_data = 8'b11111111;
		20'b00010100100001101111: color_data = 8'b11111111;
		20'b00010100100001110000: color_data = 8'b11111111;
		20'b00010100100001110001: color_data = 8'b11111111;
		20'b00010100100001110010: color_data = 8'b11111111;
		20'b00010100100001110011: color_data = 8'b11111111;
		20'b00010100100001110100: color_data = 8'b11111111;
		20'b00010100100001110101: color_data = 8'b11111111;
		20'b00010100100001110110: color_data = 8'b11111111;
		20'b00010100100001110111: color_data = 8'b11111111;
		20'b00010100100001111000: color_data = 8'b11111111;
		20'b00010100100001111001: color_data = 8'b11111111;
		20'b00010100100001111010: color_data = 8'b11111111;
		20'b00010100100001111011: color_data = 8'b11111111;
		20'b00010100100001111100: color_data = 8'b11111111;
		20'b00010100100001111101: color_data = 8'b11111111;
		20'b00010100100001111110: color_data = 8'b11111111;
		20'b00010100100001111111: color_data = 8'b11111111;
		20'b00010100100010000000: color_data = 8'b11111111;
		20'b00010100100010000001: color_data = 8'b11111111;
		20'b00010100100010000010: color_data = 8'b11111111;
		20'b00010100100010000011: color_data = 8'b11111111;
		20'b00010100100010000100: color_data = 8'b11111111;
		20'b00010100100010000101: color_data = 8'b11111111;
		20'b00010100100010000110: color_data = 8'b11111111;
		20'b00010100100010000111: color_data = 8'b11111111;
		20'b00010100100010001000: color_data = 8'b11111111;
		20'b00010100100010001001: color_data = 8'b11111111;
		20'b00010100100010001010: color_data = 8'b11111111;
		20'b00010100100010001011: color_data = 8'b11111111;
		20'b00010100100010001100: color_data = 8'b11111111;
		20'b00010100100010001101: color_data = 8'b11111111;
		20'b00010100100010001110: color_data = 8'b11111111;
		20'b00010100100010011000: color_data = 8'b11011011;
		20'b00010100100010011001: color_data = 8'b11111111;
		20'b00010100100010011010: color_data = 8'b11111111;
		20'b00010100100010011011: color_data = 8'b11111111;
		20'b00010100100010011100: color_data = 8'b11111111;
		20'b00010100100010011101: color_data = 8'b11111111;
		20'b00010100100010011110: color_data = 8'b11111111;
		20'b00010100100010011111: color_data = 8'b11111111;
		20'b00010100100010100000: color_data = 8'b11111111;
		20'b00010100100010100001: color_data = 8'b11111111;
		20'b00010100100010100010: color_data = 8'b11111111;
		20'b00010100100010100011: color_data = 8'b11111111;
		20'b00010100100010100100: color_data = 8'b11111111;
		20'b00010100100010100101: color_data = 8'b11111111;
		20'b00010100100010100110: color_data = 8'b11111111;
		20'b00010100100010100111: color_data = 8'b11111111;
		20'b00010100100010101000: color_data = 8'b11111111;
		20'b00010100100010101001: color_data = 8'b11111111;
		20'b00010100100010101010: color_data = 8'b11111111;
		20'b00010100100010101011: color_data = 8'b11111111;
		20'b00010100100010101100: color_data = 8'b11111111;
		20'b00010100100010101101: color_data = 8'b11111111;
		20'b00010100100010101110: color_data = 8'b11111111;
		20'b00010100100010101111: color_data = 8'b11111111;
		20'b00010100100010110000: color_data = 8'b11111111;
		20'b00010100100010110001: color_data = 8'b11111111;
		20'b00010100100010110010: color_data = 8'b11111111;
		20'b00010100100010110011: color_data = 8'b11111111;
		20'b00010100100010110100: color_data = 8'b11111111;
		20'b00010100100010110101: color_data = 8'b11111111;
		20'b00010100100010110110: color_data = 8'b11111111;
		20'b00010100100010110111: color_data = 8'b11111111;
		20'b00010100100010111000: color_data = 8'b11111111;
		20'b00010100100010111001: color_data = 8'b11111111;
		20'b00010100100010111010: color_data = 8'b11111111;
		20'b00010100100010111011: color_data = 8'b11111111;
		20'b00010100100010111100: color_data = 8'b11111111;
		20'b00010100100010111101: color_data = 8'b11111111;
		20'b00010100100010111110: color_data = 8'b11011011;

		20'b00010100110000001001: color_data = 8'b11011011;
		20'b00010100110000001010: color_data = 8'b11111111;
		20'b00010100110000001011: color_data = 8'b11111111;
		20'b00010100110000001100: color_data = 8'b11111111;
		20'b00010100110000001101: color_data = 8'b11111111;
		20'b00010100110000001110: color_data = 8'b11111111;
		20'b00010100110000001111: color_data = 8'b11111111;
		20'b00010100110000010000: color_data = 8'b11111111;
		20'b00010100110000010001: color_data = 8'b11111111;
		20'b00010100110000010010: color_data = 8'b11111111;
		20'b00010100110000010011: color_data = 8'b11111111;
		20'b00010100110000010100: color_data = 8'b11111111;
		20'b00010100110000010101: color_data = 8'b11111111;
		20'b00010100110000010110: color_data = 8'b11111111;
		20'b00010100110000010111: color_data = 8'b11111111;
		20'b00010100110000011000: color_data = 8'b11111111;
		20'b00010100110000011001: color_data = 8'b11111111;
		20'b00010100110000011010: color_data = 8'b11111111;
		20'b00010100110000011011: color_data = 8'b11111111;
		20'b00010100110000011100: color_data = 8'b11111111;
		20'b00010100110000011101: color_data = 8'b11111111;
		20'b00010100110000011110: color_data = 8'b11111111;
		20'b00010100110000011111: color_data = 8'b11111111;
		20'b00010100110000100000: color_data = 8'b11111111;
		20'b00010100110000100001: color_data = 8'b11111111;
		20'b00010100110000100010: color_data = 8'b11111111;
		20'b00010100110000100011: color_data = 8'b11111111;
		20'b00010100110000100100: color_data = 8'b11111111;
		20'b00010100110000100101: color_data = 8'b11111111;
		20'b00010100110000100110: color_data = 8'b11111111;
		20'b00010100110000100111: color_data = 8'b11111111;
		20'b00010100110000101000: color_data = 8'b11111111;
		20'b00010100110000101001: color_data = 8'b11111111;
		20'b00010100110000101010: color_data = 8'b11111111;
		20'b00010100110000101011: color_data = 8'b11111111;
		20'b00010100110000101100: color_data = 8'b11111111;
		20'b00010100110000101101: color_data = 8'b11111111;
		20'b00010100110000101110: color_data = 8'b11111111;
		20'b00010100110000101111: color_data = 8'b11011011;
		20'b00010100110000111001: color_data = 8'b11111111;
		20'b00010100110000111010: color_data = 8'b11111111;
		20'b00010100110000111011: color_data = 8'b11111111;
		20'b00010100110000111100: color_data = 8'b11111111;
		20'b00010100110000111101: color_data = 8'b11111111;
		20'b00010100110000111110: color_data = 8'b11111111;
		20'b00010100110000111111: color_data = 8'b11111111;
		20'b00010100110001000000: color_data = 8'b11111111;
		20'b00010100110001000001: color_data = 8'b11111111;
		20'b00010100110001000010: color_data = 8'b11111111;
		20'b00010100110001000011: color_data = 8'b11111111;
		20'b00010100110001000100: color_data = 8'b11111111;
		20'b00010100110001000101: color_data = 8'b11111111;
		20'b00010100110001000110: color_data = 8'b11111111;
		20'b00010100110001000111: color_data = 8'b11111111;
		20'b00010100110001001000: color_data = 8'b11111111;
		20'b00010100110001001001: color_data = 8'b11111111;
		20'b00010100110001001010: color_data = 8'b11111111;
		20'b00010100110001001011: color_data = 8'b11111111;
		20'b00010100110001001100: color_data = 8'b11111111;
		20'b00010100110001001101: color_data = 8'b11111111;
		20'b00010100110001001110: color_data = 8'b11111111;
		20'b00010100110001001111: color_data = 8'b11111111;
		20'b00010100110001010000: color_data = 8'b11111111;
		20'b00010100110001010001: color_data = 8'b11111111;
		20'b00010100110001010010: color_data = 8'b11111111;
		20'b00010100110001010011: color_data = 8'b11111111;
		20'b00010100110001010100: color_data = 8'b11111111;
		20'b00010100110001010101: color_data = 8'b11111111;
		20'b00010100110001010110: color_data = 8'b11111111;
		20'b00010100110001010111: color_data = 8'b11111111;
		20'b00010100110001011000: color_data = 8'b11111111;
		20'b00010100110001011001: color_data = 8'b11111111;
		20'b00010100110001011010: color_data = 8'b11111111;
		20'b00010100110001011011: color_data = 8'b11111111;
		20'b00010100110001011100: color_data = 8'b11111111;
		20'b00010100110001011101: color_data = 8'b11111111;
		20'b00010100110001011110: color_data = 8'b11111111;
		20'b00010100110001011111: color_data = 8'b10010010;
		20'b00010100110001101000: color_data = 8'b10010010;
		20'b00010100110001101001: color_data = 8'b11111111;
		20'b00010100110001101010: color_data = 8'b11111111;
		20'b00010100110001101011: color_data = 8'b11111111;
		20'b00010100110001101100: color_data = 8'b11111111;
		20'b00010100110001101101: color_data = 8'b11111111;
		20'b00010100110001101110: color_data = 8'b11111111;
		20'b00010100110001101111: color_data = 8'b11111111;
		20'b00010100110001110000: color_data = 8'b11111111;
		20'b00010100110001110001: color_data = 8'b11111111;
		20'b00010100110001110010: color_data = 8'b11111111;
		20'b00010100110001110011: color_data = 8'b11111111;
		20'b00010100110001110100: color_data = 8'b11111111;
		20'b00010100110001110101: color_data = 8'b11111111;
		20'b00010100110001110110: color_data = 8'b11111111;
		20'b00010100110001110111: color_data = 8'b11111111;
		20'b00010100110001111000: color_data = 8'b11111111;
		20'b00010100110001111001: color_data = 8'b11111111;
		20'b00010100110001111010: color_data = 8'b11111111;
		20'b00010100110001111011: color_data = 8'b11111111;
		20'b00010100110001111100: color_data = 8'b11111111;
		20'b00010100110001111101: color_data = 8'b11111111;
		20'b00010100110001111110: color_data = 8'b11111111;
		20'b00010100110001111111: color_data = 8'b11111111;
		20'b00010100110010000000: color_data = 8'b11111111;
		20'b00010100110010000001: color_data = 8'b11111111;
		20'b00010100110010000010: color_data = 8'b11111111;
		20'b00010100110010000011: color_data = 8'b11111111;
		20'b00010100110010000100: color_data = 8'b11111111;
		20'b00010100110010000101: color_data = 8'b11111111;
		20'b00010100110010000110: color_data = 8'b11111111;
		20'b00010100110010000111: color_data = 8'b11111111;
		20'b00010100110010001000: color_data = 8'b11111111;
		20'b00010100110010001001: color_data = 8'b11111111;
		20'b00010100110010001010: color_data = 8'b11111111;
		20'b00010100110010001011: color_data = 8'b11111111;
		20'b00010100110010001100: color_data = 8'b11111111;
		20'b00010100110010001101: color_data = 8'b11111111;
		20'b00010100110010001110: color_data = 8'b11111111;
		20'b00010100110010011000: color_data = 8'b11011011;
		20'b00010100110010011001: color_data = 8'b11111111;
		20'b00010100110010011010: color_data = 8'b11111111;
		20'b00010100110010011011: color_data = 8'b11111111;
		20'b00010100110010011100: color_data = 8'b11111111;
		20'b00010100110010011101: color_data = 8'b11111111;
		20'b00010100110010011110: color_data = 8'b11111111;
		20'b00010100110010011111: color_data = 8'b11111111;
		20'b00010100110010100000: color_data = 8'b11111111;
		20'b00010100110010100001: color_data = 8'b11111111;
		20'b00010100110010100010: color_data = 8'b11111111;
		20'b00010100110010100011: color_data = 8'b11111111;
		20'b00010100110010100100: color_data = 8'b11111111;
		20'b00010100110010100101: color_data = 8'b11111111;
		20'b00010100110010100110: color_data = 8'b11111111;
		20'b00010100110010100111: color_data = 8'b11111111;
		20'b00010100110010101000: color_data = 8'b11111111;
		20'b00010100110010101001: color_data = 8'b11111111;
		20'b00010100110010101010: color_data = 8'b11111111;
		20'b00010100110010101011: color_data = 8'b11111111;
		20'b00010100110010101100: color_data = 8'b11111111;
		20'b00010100110010101101: color_data = 8'b11111111;
		20'b00010100110010101110: color_data = 8'b11111111;
		20'b00010100110010101111: color_data = 8'b11111111;
		20'b00010100110010110000: color_data = 8'b11111111;
		20'b00010100110010110001: color_data = 8'b11111111;
		20'b00010100110010110010: color_data = 8'b11111111;
		20'b00010100110010110011: color_data = 8'b11111111;
		20'b00010100110010110100: color_data = 8'b11111111;
		20'b00010100110010110101: color_data = 8'b11111111;
		20'b00010100110010110110: color_data = 8'b11111111;
		20'b00010100110010110111: color_data = 8'b11111111;
		20'b00010100110010111000: color_data = 8'b11111111;
		20'b00010100110010111001: color_data = 8'b11111111;
		20'b00010100110010111010: color_data = 8'b11111111;
		20'b00010100110010111011: color_data = 8'b11111111;
		20'b00010100110010111100: color_data = 8'b11111111;
		20'b00010100110010111101: color_data = 8'b11111111;
		20'b00010100110010111110: color_data = 8'b11011011;

		20'b00010101000000001001: color_data = 8'b11011011;
		20'b00010101000000001010: color_data = 8'b11111111;
		20'b00010101000000001011: color_data = 8'b11111111;
		20'b00010101000000001100: color_data = 8'b11111111;
		20'b00010101000000001101: color_data = 8'b11111111;
		20'b00010101000000001110: color_data = 8'b11111111;
		20'b00010101000000001111: color_data = 8'b11111111;
		20'b00010101000000010000: color_data = 8'b11111111;
		20'b00010101000000010001: color_data = 8'b11111111;
		20'b00010101000000010010: color_data = 8'b11111111;
		20'b00010101000000010011: color_data = 8'b11111111;
		20'b00010101000000010100: color_data = 8'b11111111;
		20'b00010101000000010101: color_data = 8'b11111111;
		20'b00010101000000010110: color_data = 8'b11111111;
		20'b00010101000000010111: color_data = 8'b11111111;
		20'b00010101000000011000: color_data = 8'b11111111;
		20'b00010101000000011001: color_data = 8'b11111111;
		20'b00010101000000011010: color_data = 8'b11111111;
		20'b00010101000000011011: color_data = 8'b11111111;
		20'b00010101000000011100: color_data = 8'b11111111;
		20'b00010101000000011101: color_data = 8'b11111111;
		20'b00010101000000011110: color_data = 8'b11111111;
		20'b00010101000000011111: color_data = 8'b11111111;
		20'b00010101000000100000: color_data = 8'b11111111;
		20'b00010101000000100001: color_data = 8'b11111111;
		20'b00010101000000100010: color_data = 8'b11111111;
		20'b00010101000000100011: color_data = 8'b11111111;
		20'b00010101000000100100: color_data = 8'b11111111;
		20'b00010101000000100101: color_data = 8'b11111111;
		20'b00010101000000100110: color_data = 8'b11111111;
		20'b00010101000000100111: color_data = 8'b11111111;
		20'b00010101000000101000: color_data = 8'b11111111;
		20'b00010101000000101001: color_data = 8'b11111111;
		20'b00010101000000101010: color_data = 8'b11111111;
		20'b00010101000000101011: color_data = 8'b11111111;
		20'b00010101000000101100: color_data = 8'b11111111;
		20'b00010101000000101101: color_data = 8'b11111111;
		20'b00010101000000101110: color_data = 8'b11111111;
		20'b00010101000000101111: color_data = 8'b11011011;
		20'b00010101000000111001: color_data = 8'b11111111;
		20'b00010101000000111010: color_data = 8'b11111111;
		20'b00010101000000111011: color_data = 8'b11111111;
		20'b00010101000000111100: color_data = 8'b11111111;
		20'b00010101000000111101: color_data = 8'b11111111;
		20'b00010101000000111110: color_data = 8'b11111111;
		20'b00010101000000111111: color_data = 8'b11111111;
		20'b00010101000001000000: color_data = 8'b11111111;
		20'b00010101000001000001: color_data = 8'b11111111;
		20'b00010101000001000010: color_data = 8'b11111111;
		20'b00010101000001000011: color_data = 8'b11111111;
		20'b00010101000001000100: color_data = 8'b11111111;
		20'b00010101000001000101: color_data = 8'b11111111;
		20'b00010101000001000110: color_data = 8'b11111111;
		20'b00010101000001000111: color_data = 8'b11111111;
		20'b00010101000001001000: color_data = 8'b11111111;
		20'b00010101000001001001: color_data = 8'b11111111;
		20'b00010101000001001010: color_data = 8'b11111111;
		20'b00010101000001001011: color_data = 8'b11111111;
		20'b00010101000001001100: color_data = 8'b11111111;
		20'b00010101000001001101: color_data = 8'b11111111;
		20'b00010101000001001110: color_data = 8'b11111111;
		20'b00010101000001001111: color_data = 8'b11111111;
		20'b00010101000001010000: color_data = 8'b11111111;
		20'b00010101000001010001: color_data = 8'b11111111;
		20'b00010101000001010010: color_data = 8'b11111111;
		20'b00010101000001010011: color_data = 8'b11111111;
		20'b00010101000001010100: color_data = 8'b11111111;
		20'b00010101000001010101: color_data = 8'b11111111;
		20'b00010101000001010110: color_data = 8'b11111111;
		20'b00010101000001010111: color_data = 8'b11111111;
		20'b00010101000001011000: color_data = 8'b11111111;
		20'b00010101000001011001: color_data = 8'b11111111;
		20'b00010101000001011010: color_data = 8'b11111111;
		20'b00010101000001011011: color_data = 8'b11111111;
		20'b00010101000001011100: color_data = 8'b11111111;
		20'b00010101000001011101: color_data = 8'b11111111;
		20'b00010101000001011110: color_data = 8'b11111111;
		20'b00010101000001011111: color_data = 8'b10010010;
		20'b00010101000001101000: color_data = 8'b10010010;
		20'b00010101000001101001: color_data = 8'b11111111;
		20'b00010101000001101010: color_data = 8'b11111111;
		20'b00010101000001101011: color_data = 8'b11111111;
		20'b00010101000001101100: color_data = 8'b11111111;
		20'b00010101000001101101: color_data = 8'b11111111;
		20'b00010101000001101110: color_data = 8'b11111111;
		20'b00010101000001101111: color_data = 8'b11111111;
		20'b00010101000001110000: color_data = 8'b11111111;
		20'b00010101000001110001: color_data = 8'b11111111;
		20'b00010101000001110010: color_data = 8'b11111111;
		20'b00010101000001110011: color_data = 8'b11111111;
		20'b00010101000001110100: color_data = 8'b11111111;
		20'b00010101000001110101: color_data = 8'b11111111;
		20'b00010101000001110110: color_data = 8'b11111111;
		20'b00010101000001110111: color_data = 8'b11111111;
		20'b00010101000001111000: color_data = 8'b11111111;
		20'b00010101000001111001: color_data = 8'b11111111;
		20'b00010101000001111010: color_data = 8'b11111111;
		20'b00010101000001111011: color_data = 8'b11111111;
		20'b00010101000001111100: color_data = 8'b11111111;
		20'b00010101000001111101: color_data = 8'b11111111;
		20'b00010101000001111110: color_data = 8'b11111111;
		20'b00010101000001111111: color_data = 8'b11111111;
		20'b00010101000010000000: color_data = 8'b11111111;
		20'b00010101000010000001: color_data = 8'b11111111;
		20'b00010101000010000010: color_data = 8'b11111111;
		20'b00010101000010000011: color_data = 8'b11111111;
		20'b00010101000010000100: color_data = 8'b11111111;
		20'b00010101000010000101: color_data = 8'b11111111;
		20'b00010101000010000110: color_data = 8'b11111111;
		20'b00010101000010000111: color_data = 8'b11111111;
		20'b00010101000010001000: color_data = 8'b11111111;
		20'b00010101000010001001: color_data = 8'b11111111;
		20'b00010101000010001010: color_data = 8'b11111111;
		20'b00010101000010001011: color_data = 8'b11111111;
		20'b00010101000010001100: color_data = 8'b11111111;
		20'b00010101000010001101: color_data = 8'b11111111;
		20'b00010101000010001110: color_data = 8'b11111111;
		20'b00010101000010011000: color_data = 8'b11011011;
		20'b00010101000010011001: color_data = 8'b11111111;
		20'b00010101000010011010: color_data = 8'b11111111;
		20'b00010101000010011011: color_data = 8'b11111111;
		20'b00010101000010011100: color_data = 8'b11111111;
		20'b00010101000010011101: color_data = 8'b11111111;
		20'b00010101000010011110: color_data = 8'b11111111;
		20'b00010101000010011111: color_data = 8'b11111111;
		20'b00010101000010100000: color_data = 8'b11111111;
		20'b00010101000010100001: color_data = 8'b11111111;
		20'b00010101000010100010: color_data = 8'b11111111;
		20'b00010101000010100011: color_data = 8'b11111111;
		20'b00010101000010100100: color_data = 8'b11111111;
		20'b00010101000010100101: color_data = 8'b11111111;
		20'b00010101000010100110: color_data = 8'b11111111;
		20'b00010101000010100111: color_data = 8'b11111111;
		20'b00010101000010101000: color_data = 8'b11111111;
		20'b00010101000010101001: color_data = 8'b11111111;
		20'b00010101000010101010: color_data = 8'b11111111;
		20'b00010101000010101011: color_data = 8'b11111111;
		20'b00010101000010101100: color_data = 8'b11111111;
		20'b00010101000010101101: color_data = 8'b11111111;
		20'b00010101000010101110: color_data = 8'b11111111;
		20'b00010101000010101111: color_data = 8'b11111111;
		20'b00010101000010110000: color_data = 8'b11111111;
		20'b00010101000010110001: color_data = 8'b11111111;
		20'b00010101000010110010: color_data = 8'b11111111;
		20'b00010101000010110011: color_data = 8'b11111111;
		20'b00010101000010110100: color_data = 8'b11111111;
		20'b00010101000010110101: color_data = 8'b11111111;
		20'b00010101000010110110: color_data = 8'b11111111;
		20'b00010101000010110111: color_data = 8'b11111111;
		20'b00010101000010111000: color_data = 8'b11111111;
		20'b00010101000010111001: color_data = 8'b11111111;
		20'b00010101000010111010: color_data = 8'b11111111;
		20'b00010101000010111011: color_data = 8'b11111111;
		20'b00010101000010111100: color_data = 8'b11111111;
		20'b00010101000010111101: color_data = 8'b11111111;
		20'b00010101000010111110: color_data = 8'b11011011;

		20'b00010101010000001001: color_data = 8'b11011011;
		20'b00010101010000001010: color_data = 8'b11111111;
		20'b00010101010000001011: color_data = 8'b11111111;
		20'b00010101010000001100: color_data = 8'b11111111;
		20'b00010101010000001101: color_data = 8'b11111111;
		20'b00010101010000001110: color_data = 8'b11111111;
		20'b00010101010000001111: color_data = 8'b11111111;
		20'b00010101010000010000: color_data = 8'b11111111;
		20'b00010101010000010001: color_data = 8'b11111111;
		20'b00010101010000010010: color_data = 8'b11111111;
		20'b00010101010000010011: color_data = 8'b11011011;
		20'b00010101010000010100: color_data = 8'b11011011;
		20'b00010101010000010101: color_data = 8'b11011011;
		20'b00010101010000010110: color_data = 8'b11011011;
		20'b00010101010000010111: color_data = 8'b11011011;
		20'b00010101010000011000: color_data = 8'b11011011;
		20'b00010101010000011001: color_data = 8'b11011011;
		20'b00010101010000011010: color_data = 8'b11011011;
		20'b00010101010000011011: color_data = 8'b11011011;
		20'b00010101010000011100: color_data = 8'b11011011;
		20'b00010101010000011101: color_data = 8'b11011011;
		20'b00010101010000011110: color_data = 8'b11011011;
		20'b00010101010000011111: color_data = 8'b11011011;
		20'b00010101010000100000: color_data = 8'b11011011;
		20'b00010101010000100001: color_data = 8'b11011011;
		20'b00010101010000100010: color_data = 8'b11011011;
		20'b00010101010000100011: color_data = 8'b11011011;
		20'b00010101010000100100: color_data = 8'b11011011;
		20'b00010101010000100101: color_data = 8'b10010010;
		20'b00010101010000100110: color_data = 8'b11111111;
		20'b00010101010000100111: color_data = 8'b11111111;
		20'b00010101010000101000: color_data = 8'b11111111;
		20'b00010101010000101001: color_data = 8'b11111111;
		20'b00010101010000101010: color_data = 8'b11111111;
		20'b00010101010000101011: color_data = 8'b11111111;
		20'b00010101010000101100: color_data = 8'b11111111;
		20'b00010101010000101101: color_data = 8'b11111111;
		20'b00010101010000101110: color_data = 8'b11111111;
		20'b00010101010000101111: color_data = 8'b11011011;
		20'b00010101010000111001: color_data = 8'b11111111;
		20'b00010101010000111010: color_data = 8'b11111111;
		20'b00010101010000111011: color_data = 8'b11111111;
		20'b00010101010000111100: color_data = 8'b11111111;
		20'b00010101010000111101: color_data = 8'b11111111;
		20'b00010101010000111110: color_data = 8'b11111111;
		20'b00010101010000111111: color_data = 8'b11111111;
		20'b00010101010001000000: color_data = 8'b11111111;
		20'b00010101010001000001: color_data = 8'b11111111;
		20'b00010101010001000010: color_data = 8'b11111111;
		20'b00010101010001000011: color_data = 8'b11011011;
		20'b00010101010001000100: color_data = 8'b11011011;
		20'b00010101010001000101: color_data = 8'b11011011;
		20'b00010101010001000110: color_data = 8'b11011011;
		20'b00010101010001000111: color_data = 8'b11011011;
		20'b00010101010001001000: color_data = 8'b11011011;
		20'b00010101010001001001: color_data = 8'b11011011;
		20'b00010101010001001010: color_data = 8'b11011011;
		20'b00010101010001001011: color_data = 8'b11011011;
		20'b00010101010001001100: color_data = 8'b11011011;
		20'b00010101010001001101: color_data = 8'b11011011;
		20'b00010101010001001110: color_data = 8'b11011011;
		20'b00010101010001001111: color_data = 8'b11011011;
		20'b00010101010001010000: color_data = 8'b11011011;
		20'b00010101010001010001: color_data = 8'b11011011;
		20'b00010101010001010010: color_data = 8'b11011011;
		20'b00010101010001010011: color_data = 8'b11011011;
		20'b00010101010001010100: color_data = 8'b11011011;
		20'b00010101010001010101: color_data = 8'b11011011;
		20'b00010101010001010110: color_data = 8'b11111111;
		20'b00010101010001010111: color_data = 8'b11111111;
		20'b00010101010001011000: color_data = 8'b11111111;
		20'b00010101010001011001: color_data = 8'b11111111;
		20'b00010101010001011010: color_data = 8'b11111111;
		20'b00010101010001011011: color_data = 8'b11111111;
		20'b00010101010001011100: color_data = 8'b11111111;
		20'b00010101010001011101: color_data = 8'b11111111;
		20'b00010101010001011110: color_data = 8'b11111111;
		20'b00010101010001011111: color_data = 8'b10010010;
		20'b00010101010001101000: color_data = 8'b10010010;
		20'b00010101010001101001: color_data = 8'b11111111;
		20'b00010101010001101010: color_data = 8'b11111111;
		20'b00010101010001101011: color_data = 8'b11111111;
		20'b00010101010001101100: color_data = 8'b11111111;
		20'b00010101010001101101: color_data = 8'b11111111;
		20'b00010101010001101110: color_data = 8'b11111111;
		20'b00010101010001101111: color_data = 8'b11111111;
		20'b00010101010001110000: color_data = 8'b11111111;
		20'b00010101010001110001: color_data = 8'b11111111;
		20'b00010101010001110010: color_data = 8'b11011011;
		20'b00010101010001110011: color_data = 8'b11011011;
		20'b00010101010001110100: color_data = 8'b11011011;
		20'b00010101010001110101: color_data = 8'b11011011;
		20'b00010101010001110110: color_data = 8'b11011011;
		20'b00010101010001110111: color_data = 8'b11011011;
		20'b00010101010001111000: color_data = 8'b11011011;
		20'b00010101010001111001: color_data = 8'b11011011;
		20'b00010101010001111010: color_data = 8'b11011011;
		20'b00010101010001111011: color_data = 8'b11011011;
		20'b00010101010001111100: color_data = 8'b11011011;
		20'b00010101010001111101: color_data = 8'b11011011;
		20'b00010101010001111110: color_data = 8'b11011011;
		20'b00010101010001111111: color_data = 8'b11011011;
		20'b00010101010010000000: color_data = 8'b11011011;
		20'b00010101010010000001: color_data = 8'b11011011;
		20'b00010101010010000010: color_data = 8'b11011011;
		20'b00010101010010000011: color_data = 8'b11011011;
		20'b00010101010010000100: color_data = 8'b11011011;
		20'b00010101010010000101: color_data = 8'b11111111;
		20'b00010101010010000110: color_data = 8'b11111111;
		20'b00010101010010000111: color_data = 8'b11111111;
		20'b00010101010010001000: color_data = 8'b11111111;
		20'b00010101010010001001: color_data = 8'b11111111;
		20'b00010101010010001010: color_data = 8'b11111111;
		20'b00010101010010001011: color_data = 8'b11111111;
		20'b00010101010010001100: color_data = 8'b11111111;
		20'b00010101010010001101: color_data = 8'b11111111;
		20'b00010101010010001110: color_data = 8'b11111111;
		20'b00010101010010011000: color_data = 8'b11011011;
		20'b00010101010010011001: color_data = 8'b11111111;
		20'b00010101010010011010: color_data = 8'b11111111;
		20'b00010101010010011011: color_data = 8'b11111111;
		20'b00010101010010011100: color_data = 8'b11111111;
		20'b00010101010010011101: color_data = 8'b11111111;
		20'b00010101010010011110: color_data = 8'b11111111;
		20'b00010101010010011111: color_data = 8'b11111111;
		20'b00010101010010100000: color_data = 8'b11111111;
		20'b00010101010010100001: color_data = 8'b11111111;
		20'b00010101010010100010: color_data = 8'b10010010;
		20'b00010101010010100011: color_data = 8'b11011011;
		20'b00010101010010100100: color_data = 8'b11011011;
		20'b00010101010010100101: color_data = 8'b11011011;
		20'b00010101010010100110: color_data = 8'b11011011;
		20'b00010101010010100111: color_data = 8'b11011011;
		20'b00010101010010101000: color_data = 8'b11011011;
		20'b00010101010010101001: color_data = 8'b11011011;
		20'b00010101010010101010: color_data = 8'b11011011;
		20'b00010101010010101011: color_data = 8'b11011011;
		20'b00010101010010101100: color_data = 8'b11011011;
		20'b00010101010010101101: color_data = 8'b11011011;
		20'b00010101010010101110: color_data = 8'b11011011;
		20'b00010101010010101111: color_data = 8'b11011011;
		20'b00010101010010110000: color_data = 8'b11011011;
		20'b00010101010010110001: color_data = 8'b11011011;
		20'b00010101010010110010: color_data = 8'b11011011;
		20'b00010101010010110011: color_data = 8'b11011011;
		20'b00010101010010110100: color_data = 8'b11011011;
		20'b00010101010010110101: color_data = 8'b11011011;
		20'b00010101010010110110: color_data = 8'b11011011;
		20'b00010101010010110111: color_data = 8'b11011011;
		20'b00010101010010111000: color_data = 8'b11011011;
		20'b00010101010010111001: color_data = 8'b11011011;
		20'b00010101010010111010: color_data = 8'b11011011;
		20'b00010101010010111011: color_data = 8'b11011011;
		20'b00010101010010111100: color_data = 8'b11011011;
		20'b00010101010010111101: color_data = 8'b11011011;
		20'b00010101010010111110: color_data = 8'b10010010;

		20'b00010101100000001001: color_data = 8'b11011011;
		20'b00010101100000001010: color_data = 8'b11111111;
		20'b00010101100000001011: color_data = 8'b11111111;
		20'b00010101100000001100: color_data = 8'b11111111;
		20'b00010101100000001101: color_data = 8'b11111111;
		20'b00010101100000001110: color_data = 8'b11111111;
		20'b00010101100000001111: color_data = 8'b11111111;
		20'b00010101100000010000: color_data = 8'b11111111;
		20'b00010101100000010001: color_data = 8'b11111111;
		20'b00010101100000010010: color_data = 8'b11111111;
		20'b00010101100000010011: color_data = 8'b10010010;
		20'b00010101100000100110: color_data = 8'b11011011;
		20'b00010101100000100111: color_data = 8'b11111111;
		20'b00010101100000101000: color_data = 8'b11111111;
		20'b00010101100000101001: color_data = 8'b11111111;
		20'b00010101100000101010: color_data = 8'b11111111;
		20'b00010101100000101011: color_data = 8'b11111111;
		20'b00010101100000101100: color_data = 8'b11111111;
		20'b00010101100000101101: color_data = 8'b11111111;
		20'b00010101100000101110: color_data = 8'b11111111;
		20'b00010101100000101111: color_data = 8'b11011011;
		20'b00010101100000111001: color_data = 8'b11111111;
		20'b00010101100000111010: color_data = 8'b11111111;
		20'b00010101100000111011: color_data = 8'b11111111;
		20'b00010101100000111100: color_data = 8'b11111111;
		20'b00010101100000111101: color_data = 8'b11111111;
		20'b00010101100000111110: color_data = 8'b11111111;
		20'b00010101100000111111: color_data = 8'b11111111;
		20'b00010101100001000000: color_data = 8'b11111111;
		20'b00010101100001000001: color_data = 8'b11111111;
		20'b00010101100001000010: color_data = 8'b11011011;
		20'b00010101100001010101: color_data = 8'b10010010;
		20'b00010101100001010110: color_data = 8'b11111111;
		20'b00010101100001010111: color_data = 8'b11111111;
		20'b00010101100001011000: color_data = 8'b11111111;
		20'b00010101100001011001: color_data = 8'b11111111;
		20'b00010101100001011010: color_data = 8'b11111111;
		20'b00010101100001011011: color_data = 8'b11111111;
		20'b00010101100001011100: color_data = 8'b11111111;
		20'b00010101100001011101: color_data = 8'b11111111;
		20'b00010101100001011110: color_data = 8'b11111111;
		20'b00010101100001011111: color_data = 8'b10010010;
		20'b00010101100001101000: color_data = 8'b10010010;
		20'b00010101100001101001: color_data = 8'b11111111;
		20'b00010101100001101010: color_data = 8'b11111111;
		20'b00010101100001101011: color_data = 8'b11111111;
		20'b00010101100001101100: color_data = 8'b11111111;
		20'b00010101100001101101: color_data = 8'b11111111;
		20'b00010101100001101110: color_data = 8'b11111111;
		20'b00010101100001101111: color_data = 8'b11111111;
		20'b00010101100001110000: color_data = 8'b11111111;
		20'b00010101100001110001: color_data = 8'b11111111;
		20'b00010101100001110010: color_data = 8'b10010010;
		20'b00010101100010000101: color_data = 8'b11011011;
		20'b00010101100010000110: color_data = 8'b11111111;
		20'b00010101100010000111: color_data = 8'b11111111;
		20'b00010101100010001000: color_data = 8'b11111111;
		20'b00010101100010001001: color_data = 8'b11111111;
		20'b00010101100010001010: color_data = 8'b11111111;
		20'b00010101100010001011: color_data = 8'b11111111;
		20'b00010101100010001100: color_data = 8'b11111111;
		20'b00010101100010001101: color_data = 8'b11111111;
		20'b00010101100010001110: color_data = 8'b11111111;
		20'b00010101100010011000: color_data = 8'b11011011;
		20'b00010101100010011001: color_data = 8'b11111111;
		20'b00010101100010011010: color_data = 8'b11111111;
		20'b00010101100010011011: color_data = 8'b11111111;
		20'b00010101100010011100: color_data = 8'b11111111;
		20'b00010101100010011101: color_data = 8'b11111111;
		20'b00010101100010011110: color_data = 8'b11111111;
		20'b00010101100010011111: color_data = 8'b11111111;
		20'b00010101100010100000: color_data = 8'b11111111;
		20'b00010101100010100001: color_data = 8'b11011011;

		20'b00010101110000001001: color_data = 8'b11011011;
		20'b00010101110000001010: color_data = 8'b11111111;
		20'b00010101110000001011: color_data = 8'b11111111;
		20'b00010101110000001100: color_data = 8'b11111111;
		20'b00010101110000001101: color_data = 8'b11111111;
		20'b00010101110000001110: color_data = 8'b11111111;
		20'b00010101110000001111: color_data = 8'b11111111;
		20'b00010101110000010000: color_data = 8'b11111111;
		20'b00010101110000010001: color_data = 8'b11111111;
		20'b00010101110000010010: color_data = 8'b11111111;
		20'b00010101110000010011: color_data = 8'b10010010;
		20'b00010101110000100110: color_data = 8'b11011011;
		20'b00010101110000100111: color_data = 8'b11111111;
		20'b00010101110000101000: color_data = 8'b11111111;
		20'b00010101110000101001: color_data = 8'b11111111;
		20'b00010101110000101010: color_data = 8'b11111111;
		20'b00010101110000101011: color_data = 8'b11111111;
		20'b00010101110000101100: color_data = 8'b11111111;
		20'b00010101110000101101: color_data = 8'b11111111;
		20'b00010101110000101110: color_data = 8'b11111111;
		20'b00010101110000101111: color_data = 8'b11011011;
		20'b00010101110000111001: color_data = 8'b11111111;
		20'b00010101110000111010: color_data = 8'b11111111;
		20'b00010101110000111011: color_data = 8'b11111111;
		20'b00010101110000111100: color_data = 8'b11111111;
		20'b00010101110000111101: color_data = 8'b11111111;
		20'b00010101110000111110: color_data = 8'b11111111;
		20'b00010101110000111111: color_data = 8'b11111111;
		20'b00010101110001000000: color_data = 8'b11111111;
		20'b00010101110001000001: color_data = 8'b11111111;
		20'b00010101110001000010: color_data = 8'b11011011;
		20'b00010101110001010101: color_data = 8'b10010010;
		20'b00010101110001010110: color_data = 8'b11111111;
		20'b00010101110001010111: color_data = 8'b11111111;
		20'b00010101110001011000: color_data = 8'b11111111;
		20'b00010101110001011001: color_data = 8'b11111111;
		20'b00010101110001011010: color_data = 8'b11111111;
		20'b00010101110001011011: color_data = 8'b11111111;
		20'b00010101110001011100: color_data = 8'b11111111;
		20'b00010101110001011101: color_data = 8'b11111111;
		20'b00010101110001011110: color_data = 8'b11111111;
		20'b00010101110001011111: color_data = 8'b10010010;
		20'b00010101110001101000: color_data = 8'b10010010;
		20'b00010101110001101001: color_data = 8'b11111111;
		20'b00010101110001101010: color_data = 8'b11111111;
		20'b00010101110001101011: color_data = 8'b11111111;
		20'b00010101110001101100: color_data = 8'b11111111;
		20'b00010101110001101101: color_data = 8'b11111111;
		20'b00010101110001101110: color_data = 8'b11111111;
		20'b00010101110001101111: color_data = 8'b11111111;
		20'b00010101110001110000: color_data = 8'b11111111;
		20'b00010101110001110001: color_data = 8'b11111111;
		20'b00010101110001110010: color_data = 8'b10010010;
		20'b00010101110010000101: color_data = 8'b11011011;
		20'b00010101110010000110: color_data = 8'b11111111;
		20'b00010101110010000111: color_data = 8'b11111111;
		20'b00010101110010001000: color_data = 8'b11111111;
		20'b00010101110010001001: color_data = 8'b11111111;
		20'b00010101110010001010: color_data = 8'b11111111;
		20'b00010101110010001011: color_data = 8'b11111111;
		20'b00010101110010001100: color_data = 8'b11111111;
		20'b00010101110010001101: color_data = 8'b11111111;
		20'b00010101110010001110: color_data = 8'b11111111;
		20'b00010101110010011000: color_data = 8'b11011011;
		20'b00010101110010011001: color_data = 8'b11111111;
		20'b00010101110010011010: color_data = 8'b11111111;
		20'b00010101110010011011: color_data = 8'b11111111;
		20'b00010101110010011100: color_data = 8'b11111111;
		20'b00010101110010011101: color_data = 8'b11111111;
		20'b00010101110010011110: color_data = 8'b11111111;
		20'b00010101110010011111: color_data = 8'b11111111;
		20'b00010101110010100000: color_data = 8'b11111111;
		20'b00010101110010100001: color_data = 8'b11011011;

		20'b00010110000000001001: color_data = 8'b11011011;
		20'b00010110000000001010: color_data = 8'b11111111;
		20'b00010110000000001011: color_data = 8'b11111111;
		20'b00010110000000001100: color_data = 8'b11111111;
		20'b00010110000000001101: color_data = 8'b11111111;
		20'b00010110000000001110: color_data = 8'b11111111;
		20'b00010110000000001111: color_data = 8'b11111111;
		20'b00010110000000010000: color_data = 8'b11111111;
		20'b00010110000000010001: color_data = 8'b11111111;
		20'b00010110000000010010: color_data = 8'b11111111;
		20'b00010110000000010011: color_data = 8'b10010010;
		20'b00010110000000100110: color_data = 8'b11011011;
		20'b00010110000000100111: color_data = 8'b11111111;
		20'b00010110000000101000: color_data = 8'b11111111;
		20'b00010110000000101001: color_data = 8'b11111111;
		20'b00010110000000101010: color_data = 8'b11111111;
		20'b00010110000000101011: color_data = 8'b11111111;
		20'b00010110000000101100: color_data = 8'b11111111;
		20'b00010110000000101101: color_data = 8'b11111111;
		20'b00010110000000101110: color_data = 8'b11111111;
		20'b00010110000000101111: color_data = 8'b11011011;
		20'b00010110000000111001: color_data = 8'b11111111;
		20'b00010110000000111010: color_data = 8'b11111111;
		20'b00010110000000111011: color_data = 8'b11111111;
		20'b00010110000000111100: color_data = 8'b11111111;
		20'b00010110000000111101: color_data = 8'b11111111;
		20'b00010110000000111110: color_data = 8'b11111111;
		20'b00010110000000111111: color_data = 8'b11111111;
		20'b00010110000001000000: color_data = 8'b11111111;
		20'b00010110000001000001: color_data = 8'b11111111;
		20'b00010110000001000010: color_data = 8'b11011011;
		20'b00010110000001010101: color_data = 8'b10010010;
		20'b00010110000001010110: color_data = 8'b11111111;
		20'b00010110000001010111: color_data = 8'b11111111;
		20'b00010110000001011000: color_data = 8'b11111111;
		20'b00010110000001011001: color_data = 8'b11111111;
		20'b00010110000001011010: color_data = 8'b11111111;
		20'b00010110000001011011: color_data = 8'b11111111;
		20'b00010110000001011100: color_data = 8'b11111111;
		20'b00010110000001011101: color_data = 8'b11111111;
		20'b00010110000001011110: color_data = 8'b11111111;
		20'b00010110000001011111: color_data = 8'b10010010;
		20'b00010110000001101000: color_data = 8'b10010010;
		20'b00010110000001101001: color_data = 8'b11111111;
		20'b00010110000001101010: color_data = 8'b11111111;
		20'b00010110000001101011: color_data = 8'b11111111;
		20'b00010110000001101100: color_data = 8'b11111111;
		20'b00010110000001101101: color_data = 8'b11111111;
		20'b00010110000001101110: color_data = 8'b11111111;
		20'b00010110000001101111: color_data = 8'b11111111;
		20'b00010110000001110000: color_data = 8'b11111111;
		20'b00010110000001110001: color_data = 8'b11111111;
		20'b00010110000001110010: color_data = 8'b10010010;
		20'b00010110000010000101: color_data = 8'b11011011;
		20'b00010110000010000110: color_data = 8'b11111111;
		20'b00010110000010000111: color_data = 8'b11111111;
		20'b00010110000010001000: color_data = 8'b11111111;
		20'b00010110000010001001: color_data = 8'b11111111;
		20'b00010110000010001010: color_data = 8'b11111111;
		20'b00010110000010001011: color_data = 8'b11111111;
		20'b00010110000010001100: color_data = 8'b11111111;
		20'b00010110000010001101: color_data = 8'b11111111;
		20'b00010110000010001110: color_data = 8'b11111111;
		20'b00010110000010011000: color_data = 8'b11011011;
		20'b00010110000010011001: color_data = 8'b11111111;
		20'b00010110000010011010: color_data = 8'b11111111;
		20'b00010110000010011011: color_data = 8'b11111111;
		20'b00010110000010011100: color_data = 8'b11111111;
		20'b00010110000010011101: color_data = 8'b11111111;
		20'b00010110000010011110: color_data = 8'b11111111;
		20'b00010110000010011111: color_data = 8'b11111111;
		20'b00010110000010100000: color_data = 8'b11111111;
		20'b00010110000010100001: color_data = 8'b11011011;

		20'b00010110010000001001: color_data = 8'b11011011;
		20'b00010110010000001010: color_data = 8'b11111111;
		20'b00010110010000001011: color_data = 8'b11111111;
		20'b00010110010000001100: color_data = 8'b11111111;
		20'b00010110010000001101: color_data = 8'b11111111;
		20'b00010110010000001110: color_data = 8'b11111111;
		20'b00010110010000001111: color_data = 8'b11111111;
		20'b00010110010000010000: color_data = 8'b11111111;
		20'b00010110010000010001: color_data = 8'b11111111;
		20'b00010110010000010010: color_data = 8'b11111111;
		20'b00010110010000010011: color_data = 8'b10010010;
		20'b00010110010000100110: color_data = 8'b11011011;
		20'b00010110010000100111: color_data = 8'b11111111;
		20'b00010110010000101000: color_data = 8'b11111111;
		20'b00010110010000101001: color_data = 8'b11111111;
		20'b00010110010000101010: color_data = 8'b11111111;
		20'b00010110010000101011: color_data = 8'b11111111;
		20'b00010110010000101100: color_data = 8'b11111111;
		20'b00010110010000101101: color_data = 8'b11111111;
		20'b00010110010000101110: color_data = 8'b11111111;
		20'b00010110010000101111: color_data = 8'b11011011;
		20'b00010110010000111001: color_data = 8'b11111111;
		20'b00010110010000111010: color_data = 8'b11111111;
		20'b00010110010000111011: color_data = 8'b11111111;
		20'b00010110010000111100: color_data = 8'b11111111;
		20'b00010110010000111101: color_data = 8'b11111111;
		20'b00010110010000111110: color_data = 8'b11111111;
		20'b00010110010000111111: color_data = 8'b11111111;
		20'b00010110010001000000: color_data = 8'b11111111;
		20'b00010110010001000001: color_data = 8'b11111111;
		20'b00010110010001000010: color_data = 8'b11011011;
		20'b00010110010001010101: color_data = 8'b10010010;
		20'b00010110010001010110: color_data = 8'b11111111;
		20'b00010110010001010111: color_data = 8'b11111111;
		20'b00010110010001011000: color_data = 8'b11111111;
		20'b00010110010001011001: color_data = 8'b11111111;
		20'b00010110010001011010: color_data = 8'b11111111;
		20'b00010110010001011011: color_data = 8'b11111111;
		20'b00010110010001011100: color_data = 8'b11111111;
		20'b00010110010001011101: color_data = 8'b11111111;
		20'b00010110010001011110: color_data = 8'b11111111;
		20'b00010110010001011111: color_data = 8'b10010010;
		20'b00010110010001101000: color_data = 8'b10010010;
		20'b00010110010001101001: color_data = 8'b11111111;
		20'b00010110010001101010: color_data = 8'b11111111;
		20'b00010110010001101011: color_data = 8'b11111111;
		20'b00010110010001101100: color_data = 8'b11111111;
		20'b00010110010001101101: color_data = 8'b11111111;
		20'b00010110010001101110: color_data = 8'b11111111;
		20'b00010110010001101111: color_data = 8'b11111111;
		20'b00010110010001110000: color_data = 8'b11111111;
		20'b00010110010001110001: color_data = 8'b11111111;
		20'b00010110010001110010: color_data = 8'b10010010;
		20'b00010110010010000101: color_data = 8'b11011011;
		20'b00010110010010000110: color_data = 8'b11111111;
		20'b00010110010010000111: color_data = 8'b11111111;
		20'b00010110010010001000: color_data = 8'b11111111;
		20'b00010110010010001001: color_data = 8'b11111111;
		20'b00010110010010001010: color_data = 8'b11111111;
		20'b00010110010010001011: color_data = 8'b11111111;
		20'b00010110010010001100: color_data = 8'b11111111;
		20'b00010110010010001101: color_data = 8'b11111111;
		20'b00010110010010001110: color_data = 8'b11111111;
		20'b00010110010010011000: color_data = 8'b11011011;
		20'b00010110010010011001: color_data = 8'b11111111;
		20'b00010110010010011010: color_data = 8'b11111111;
		20'b00010110010010011011: color_data = 8'b11111111;
		20'b00010110010010011100: color_data = 8'b11111111;
		20'b00010110010010011101: color_data = 8'b11111111;
		20'b00010110010010011110: color_data = 8'b11111111;
		20'b00010110010010011111: color_data = 8'b11111111;
		20'b00010110010010100000: color_data = 8'b11111111;
		20'b00010110010010100001: color_data = 8'b11011011;

		20'b00010110100000001001: color_data = 8'b11011011;
		20'b00010110100000001010: color_data = 8'b11111111;
		20'b00010110100000001011: color_data = 8'b11111111;
		20'b00010110100000001100: color_data = 8'b11111111;
		20'b00010110100000001101: color_data = 8'b11111111;
		20'b00010110100000001110: color_data = 8'b11111111;
		20'b00010110100000001111: color_data = 8'b11111111;
		20'b00010110100000010000: color_data = 8'b11111111;
		20'b00010110100000010001: color_data = 8'b11111111;
		20'b00010110100000010010: color_data = 8'b11111111;
		20'b00010110100000010011: color_data = 8'b10010010;
		20'b00010110100000100110: color_data = 8'b11011011;
		20'b00010110100000100111: color_data = 8'b11111111;
		20'b00010110100000101000: color_data = 8'b11111111;
		20'b00010110100000101001: color_data = 8'b11111111;
		20'b00010110100000101010: color_data = 8'b11111111;
		20'b00010110100000101011: color_data = 8'b11111111;
		20'b00010110100000101100: color_data = 8'b11111111;
		20'b00010110100000101101: color_data = 8'b11111111;
		20'b00010110100000101110: color_data = 8'b11111111;
		20'b00010110100000101111: color_data = 8'b11011011;
		20'b00010110100000111001: color_data = 8'b11111111;
		20'b00010110100000111010: color_data = 8'b11111111;
		20'b00010110100000111011: color_data = 8'b11111111;
		20'b00010110100000111100: color_data = 8'b11111111;
		20'b00010110100000111101: color_data = 8'b11111111;
		20'b00010110100000111110: color_data = 8'b11111111;
		20'b00010110100000111111: color_data = 8'b11111111;
		20'b00010110100001000000: color_data = 8'b11111111;
		20'b00010110100001000001: color_data = 8'b11111111;
		20'b00010110100001000010: color_data = 8'b11011011;
		20'b00010110100001010101: color_data = 8'b10010010;
		20'b00010110100001010110: color_data = 8'b11111111;
		20'b00010110100001010111: color_data = 8'b11111111;
		20'b00010110100001011000: color_data = 8'b11111111;
		20'b00010110100001011001: color_data = 8'b11111111;
		20'b00010110100001011010: color_data = 8'b11111111;
		20'b00010110100001011011: color_data = 8'b11111111;
		20'b00010110100001011100: color_data = 8'b11111111;
		20'b00010110100001011101: color_data = 8'b11111111;
		20'b00010110100001011110: color_data = 8'b11111111;
		20'b00010110100001011111: color_data = 8'b10010010;
		20'b00010110100001101000: color_data = 8'b10010010;
		20'b00010110100001101001: color_data = 8'b11111111;
		20'b00010110100001101010: color_data = 8'b11111111;
		20'b00010110100001101011: color_data = 8'b11111111;
		20'b00010110100001101100: color_data = 8'b11111111;
		20'b00010110100001101101: color_data = 8'b11111111;
		20'b00010110100001101110: color_data = 8'b11111111;
		20'b00010110100001101111: color_data = 8'b11111111;
		20'b00010110100001110000: color_data = 8'b11111111;
		20'b00010110100001110001: color_data = 8'b11111111;
		20'b00010110100001110010: color_data = 8'b10010010;
		20'b00010110100010000101: color_data = 8'b11011011;
		20'b00010110100010000110: color_data = 8'b11111111;
		20'b00010110100010000111: color_data = 8'b11111111;
		20'b00010110100010001000: color_data = 8'b11111111;
		20'b00010110100010001001: color_data = 8'b11111111;
		20'b00010110100010001010: color_data = 8'b11111111;
		20'b00010110100010001011: color_data = 8'b11111111;
		20'b00010110100010001100: color_data = 8'b11111111;
		20'b00010110100010001101: color_data = 8'b11111111;
		20'b00010110100010001110: color_data = 8'b11111111;
		20'b00010110100010011000: color_data = 8'b11011011;
		20'b00010110100010011001: color_data = 8'b11111111;
		20'b00010110100010011010: color_data = 8'b11111111;
		20'b00010110100010011011: color_data = 8'b11111111;
		20'b00010110100010011100: color_data = 8'b11111111;
		20'b00010110100010011101: color_data = 8'b11111111;
		20'b00010110100010011110: color_data = 8'b11111111;
		20'b00010110100010011111: color_data = 8'b11111111;
		20'b00010110100010100000: color_data = 8'b11111111;
		20'b00010110100010100001: color_data = 8'b11011011;

		20'b00010110110000001001: color_data = 8'b11011011;
		20'b00010110110000001010: color_data = 8'b11111111;
		20'b00010110110000001011: color_data = 8'b11111111;
		20'b00010110110000001100: color_data = 8'b11111111;
		20'b00010110110000001101: color_data = 8'b11111111;
		20'b00010110110000001110: color_data = 8'b11111111;
		20'b00010110110000001111: color_data = 8'b11111111;
		20'b00010110110000010000: color_data = 8'b11111111;
		20'b00010110110000010001: color_data = 8'b11111111;
		20'b00010110110000010010: color_data = 8'b11111111;
		20'b00010110110000010011: color_data = 8'b10010010;
		20'b00010110110000100110: color_data = 8'b11011011;
		20'b00010110110000100111: color_data = 8'b11111111;
		20'b00010110110000101000: color_data = 8'b11111111;
		20'b00010110110000101001: color_data = 8'b11111111;
		20'b00010110110000101010: color_data = 8'b11111111;
		20'b00010110110000101011: color_data = 8'b11111111;
		20'b00010110110000101100: color_data = 8'b11111111;
		20'b00010110110000101101: color_data = 8'b11111111;
		20'b00010110110000101110: color_data = 8'b11111111;
		20'b00010110110000101111: color_data = 8'b11011011;
		20'b00010110110000111001: color_data = 8'b11111111;
		20'b00010110110000111010: color_data = 8'b11111111;
		20'b00010110110000111011: color_data = 8'b11111111;
		20'b00010110110000111100: color_data = 8'b11111111;
		20'b00010110110000111101: color_data = 8'b11111111;
		20'b00010110110000111110: color_data = 8'b11111111;
		20'b00010110110000111111: color_data = 8'b11111111;
		20'b00010110110001000000: color_data = 8'b11111111;
		20'b00010110110001000001: color_data = 8'b11111111;
		20'b00010110110001000010: color_data = 8'b11011011;
		20'b00010110110001010101: color_data = 8'b10010010;
		20'b00010110110001010110: color_data = 8'b11111111;
		20'b00010110110001010111: color_data = 8'b11111111;
		20'b00010110110001011000: color_data = 8'b11111111;
		20'b00010110110001011001: color_data = 8'b11111111;
		20'b00010110110001011010: color_data = 8'b11111111;
		20'b00010110110001011011: color_data = 8'b11111111;
		20'b00010110110001011100: color_data = 8'b11111111;
		20'b00010110110001011101: color_data = 8'b11111111;
		20'b00010110110001011110: color_data = 8'b11111111;
		20'b00010110110001011111: color_data = 8'b10010010;
		20'b00010110110001101000: color_data = 8'b10010010;
		20'b00010110110001101001: color_data = 8'b11111111;
		20'b00010110110001101010: color_data = 8'b11111111;
		20'b00010110110001101011: color_data = 8'b11111111;
		20'b00010110110001101100: color_data = 8'b11111111;
		20'b00010110110001101101: color_data = 8'b11111111;
		20'b00010110110001101110: color_data = 8'b11111111;
		20'b00010110110001101111: color_data = 8'b11111111;
		20'b00010110110001110000: color_data = 8'b11111111;
		20'b00010110110001110001: color_data = 8'b11111111;
		20'b00010110110001110010: color_data = 8'b10010010;
		20'b00010110110010000101: color_data = 8'b11011011;
		20'b00010110110010000110: color_data = 8'b11111111;
		20'b00010110110010000111: color_data = 8'b11111111;
		20'b00010110110010001000: color_data = 8'b11111111;
		20'b00010110110010001001: color_data = 8'b11111111;
		20'b00010110110010001010: color_data = 8'b11111111;
		20'b00010110110010001011: color_data = 8'b11111111;
		20'b00010110110010001100: color_data = 8'b11111111;
		20'b00010110110010001101: color_data = 8'b11111111;
		20'b00010110110010001110: color_data = 8'b11111111;
		20'b00010110110010011000: color_data = 8'b11011011;
		20'b00010110110010011001: color_data = 8'b11111111;
		20'b00010110110010011010: color_data = 8'b11111111;
		20'b00010110110010011011: color_data = 8'b11111111;
		20'b00010110110010011100: color_data = 8'b11111111;
		20'b00010110110010011101: color_data = 8'b11111111;
		20'b00010110110010011110: color_data = 8'b11111111;
		20'b00010110110010011111: color_data = 8'b11111111;
		20'b00010110110010100000: color_data = 8'b11111111;
		20'b00010110110010100001: color_data = 8'b11011011;

		20'b00010111000000001001: color_data = 8'b11011011;
		20'b00010111000000001010: color_data = 8'b11111111;
		20'b00010111000000001011: color_data = 8'b11111111;
		20'b00010111000000001100: color_data = 8'b11111111;
		20'b00010111000000001101: color_data = 8'b11111111;
		20'b00010111000000001110: color_data = 8'b11111111;
		20'b00010111000000001111: color_data = 8'b11111111;
		20'b00010111000000010000: color_data = 8'b11111111;
		20'b00010111000000010001: color_data = 8'b11111111;
		20'b00010111000000010010: color_data = 8'b11111111;
		20'b00010111000000010011: color_data = 8'b10010010;
		20'b00010111000000100110: color_data = 8'b11011011;
		20'b00010111000000100111: color_data = 8'b11111111;
		20'b00010111000000101000: color_data = 8'b11111111;
		20'b00010111000000101001: color_data = 8'b11111111;
		20'b00010111000000101010: color_data = 8'b11111111;
		20'b00010111000000101011: color_data = 8'b11111111;
		20'b00010111000000101100: color_data = 8'b11111111;
		20'b00010111000000101101: color_data = 8'b11111111;
		20'b00010111000000101110: color_data = 8'b11111111;
		20'b00010111000000101111: color_data = 8'b11011011;
		20'b00010111000000111001: color_data = 8'b11111111;
		20'b00010111000000111010: color_data = 8'b11111111;
		20'b00010111000000111011: color_data = 8'b11111111;
		20'b00010111000000111100: color_data = 8'b11111111;
		20'b00010111000000111101: color_data = 8'b11111111;
		20'b00010111000000111110: color_data = 8'b11111111;
		20'b00010111000000111111: color_data = 8'b11111111;
		20'b00010111000001000000: color_data = 8'b11111111;
		20'b00010111000001000001: color_data = 8'b11111111;
		20'b00010111000001000010: color_data = 8'b11011011;
		20'b00010111000001010101: color_data = 8'b10010010;
		20'b00010111000001010110: color_data = 8'b11111111;
		20'b00010111000001010111: color_data = 8'b11111111;
		20'b00010111000001011000: color_data = 8'b11111111;
		20'b00010111000001011001: color_data = 8'b11111111;
		20'b00010111000001011010: color_data = 8'b11111111;
		20'b00010111000001011011: color_data = 8'b11111111;
		20'b00010111000001011100: color_data = 8'b11111111;
		20'b00010111000001011101: color_data = 8'b11111111;
		20'b00010111000001011110: color_data = 8'b11111111;
		20'b00010111000001011111: color_data = 8'b10010010;
		20'b00010111000001101000: color_data = 8'b10010010;
		20'b00010111000001101001: color_data = 8'b11111111;
		20'b00010111000001101010: color_data = 8'b11111111;
		20'b00010111000001101011: color_data = 8'b11111111;
		20'b00010111000001101100: color_data = 8'b11111111;
		20'b00010111000001101101: color_data = 8'b11111111;
		20'b00010111000001101110: color_data = 8'b11111111;
		20'b00010111000001101111: color_data = 8'b11111111;
		20'b00010111000001110000: color_data = 8'b11111111;
		20'b00010111000001110001: color_data = 8'b11111111;
		20'b00010111000001110010: color_data = 8'b10010010;
		20'b00010111000010000101: color_data = 8'b11011011;
		20'b00010111000010000110: color_data = 8'b11111111;
		20'b00010111000010000111: color_data = 8'b11111111;
		20'b00010111000010001000: color_data = 8'b11111111;
		20'b00010111000010001001: color_data = 8'b11111111;
		20'b00010111000010001010: color_data = 8'b11111111;
		20'b00010111000010001011: color_data = 8'b11111111;
		20'b00010111000010001100: color_data = 8'b11111111;
		20'b00010111000010001101: color_data = 8'b11111111;
		20'b00010111000010001110: color_data = 8'b11111111;
		20'b00010111000010011000: color_data = 8'b11011011;
		20'b00010111000010011001: color_data = 8'b11111111;
		20'b00010111000010011010: color_data = 8'b11111111;
		20'b00010111000010011011: color_data = 8'b11111111;
		20'b00010111000010011100: color_data = 8'b11111111;
		20'b00010111000010011101: color_data = 8'b11111111;
		20'b00010111000010011110: color_data = 8'b11111111;
		20'b00010111000010011111: color_data = 8'b11111111;
		20'b00010111000010100000: color_data = 8'b11111111;
		20'b00010111000010100001: color_data = 8'b11011011;

		20'b00010111010000001001: color_data = 8'b11011011;
		20'b00010111010000001010: color_data = 8'b11111111;
		20'b00010111010000001011: color_data = 8'b11111111;
		20'b00010111010000001100: color_data = 8'b11111111;
		20'b00010111010000001101: color_data = 8'b11111111;
		20'b00010111010000001110: color_data = 8'b11111111;
		20'b00010111010000001111: color_data = 8'b11111111;
		20'b00010111010000010000: color_data = 8'b11111111;
		20'b00010111010000010001: color_data = 8'b11111111;
		20'b00010111010000010010: color_data = 8'b11111111;
		20'b00010111010000010011: color_data = 8'b10010010;
		20'b00010111010000100110: color_data = 8'b11011011;
		20'b00010111010000100111: color_data = 8'b11111111;
		20'b00010111010000101000: color_data = 8'b11111111;
		20'b00010111010000101001: color_data = 8'b11111111;
		20'b00010111010000101010: color_data = 8'b11111111;
		20'b00010111010000101011: color_data = 8'b11111111;
		20'b00010111010000101100: color_data = 8'b11111111;
		20'b00010111010000101101: color_data = 8'b11111111;
		20'b00010111010000101110: color_data = 8'b11111111;
		20'b00010111010000101111: color_data = 8'b11011011;
		20'b00010111010000111001: color_data = 8'b11111111;
		20'b00010111010000111010: color_data = 8'b11111111;
		20'b00010111010000111011: color_data = 8'b11111111;
		20'b00010111010000111100: color_data = 8'b11111111;
		20'b00010111010000111101: color_data = 8'b11111111;
		20'b00010111010000111110: color_data = 8'b11111111;
		20'b00010111010000111111: color_data = 8'b11111111;
		20'b00010111010001000000: color_data = 8'b11111111;
		20'b00010111010001000001: color_data = 8'b11111111;
		20'b00010111010001000010: color_data = 8'b11011011;
		20'b00010111010001010101: color_data = 8'b10010010;
		20'b00010111010001010110: color_data = 8'b11111111;
		20'b00010111010001010111: color_data = 8'b11111111;
		20'b00010111010001011000: color_data = 8'b11111111;
		20'b00010111010001011001: color_data = 8'b11111111;
		20'b00010111010001011010: color_data = 8'b11111111;
		20'b00010111010001011011: color_data = 8'b11111111;
		20'b00010111010001011100: color_data = 8'b11111111;
		20'b00010111010001011101: color_data = 8'b11111111;
		20'b00010111010001011110: color_data = 8'b11111111;
		20'b00010111010001011111: color_data = 8'b10010010;
		20'b00010111010001101000: color_data = 8'b10010010;
		20'b00010111010001101001: color_data = 8'b11111111;
		20'b00010111010001101010: color_data = 8'b11111111;
		20'b00010111010001101011: color_data = 8'b11111111;
		20'b00010111010001101100: color_data = 8'b11111111;
		20'b00010111010001101101: color_data = 8'b11111111;
		20'b00010111010001101110: color_data = 8'b11111111;
		20'b00010111010001101111: color_data = 8'b11111111;
		20'b00010111010001110000: color_data = 8'b11111111;
		20'b00010111010001110001: color_data = 8'b11111111;
		20'b00010111010001110010: color_data = 8'b10010010;
		20'b00010111010010000101: color_data = 8'b11011011;
		20'b00010111010010000110: color_data = 8'b11111111;
		20'b00010111010010000111: color_data = 8'b11111111;
		20'b00010111010010001000: color_data = 8'b11111111;
		20'b00010111010010001001: color_data = 8'b11111111;
		20'b00010111010010001010: color_data = 8'b11111111;
		20'b00010111010010001011: color_data = 8'b11111111;
		20'b00010111010010001100: color_data = 8'b11111111;
		20'b00010111010010001101: color_data = 8'b11111111;
		20'b00010111010010001110: color_data = 8'b11111111;
		20'b00010111010010011000: color_data = 8'b11011011;
		20'b00010111010010011001: color_data = 8'b11111111;
		20'b00010111010010011010: color_data = 8'b11111111;
		20'b00010111010010011011: color_data = 8'b11111111;
		20'b00010111010010011100: color_data = 8'b11111111;
		20'b00010111010010011101: color_data = 8'b11111111;
		20'b00010111010010011110: color_data = 8'b11111111;
		20'b00010111010010011111: color_data = 8'b11111111;
		20'b00010111010010100000: color_data = 8'b11111111;
		20'b00010111010010100001: color_data = 8'b11011011;

		20'b00010111100000001001: color_data = 8'b11011011;
		20'b00010111100000001010: color_data = 8'b11111111;
		20'b00010111100000001011: color_data = 8'b11111111;
		20'b00010111100000001100: color_data = 8'b11111111;
		20'b00010111100000001101: color_data = 8'b11111111;
		20'b00010111100000001110: color_data = 8'b11111111;
		20'b00010111100000001111: color_data = 8'b11111111;
		20'b00010111100000010000: color_data = 8'b11111111;
		20'b00010111100000010001: color_data = 8'b11111111;
		20'b00010111100000010010: color_data = 8'b11111111;
		20'b00010111100000010011: color_data = 8'b10010010;
		20'b00010111100000100110: color_data = 8'b11011011;
		20'b00010111100000100111: color_data = 8'b11111111;
		20'b00010111100000101000: color_data = 8'b11111111;
		20'b00010111100000101001: color_data = 8'b11111111;
		20'b00010111100000101010: color_data = 8'b11111111;
		20'b00010111100000101011: color_data = 8'b11111111;
		20'b00010111100000101100: color_data = 8'b11111111;
		20'b00010111100000101101: color_data = 8'b11111111;
		20'b00010111100000101110: color_data = 8'b11111111;
		20'b00010111100000101111: color_data = 8'b11011011;
		20'b00010111100000111001: color_data = 8'b11111111;
		20'b00010111100000111010: color_data = 8'b11111111;
		20'b00010111100000111011: color_data = 8'b11111111;
		20'b00010111100000111100: color_data = 8'b11111111;
		20'b00010111100000111101: color_data = 8'b11111111;
		20'b00010111100000111110: color_data = 8'b11111111;
		20'b00010111100000111111: color_data = 8'b11111111;
		20'b00010111100001000000: color_data = 8'b11111111;
		20'b00010111100001000001: color_data = 8'b11111111;
		20'b00010111100001000010: color_data = 8'b11011011;
		20'b00010111100001010101: color_data = 8'b10010010;
		20'b00010111100001010110: color_data = 8'b11111111;
		20'b00010111100001010111: color_data = 8'b11111111;
		20'b00010111100001011000: color_data = 8'b11111111;
		20'b00010111100001011001: color_data = 8'b11111111;
		20'b00010111100001011010: color_data = 8'b11111111;
		20'b00010111100001011011: color_data = 8'b11111111;
		20'b00010111100001011100: color_data = 8'b11111111;
		20'b00010111100001011101: color_data = 8'b11111111;
		20'b00010111100001011110: color_data = 8'b11111111;
		20'b00010111100001011111: color_data = 8'b10010010;
		20'b00010111100001101000: color_data = 8'b10010010;
		20'b00010111100001101001: color_data = 8'b11111111;
		20'b00010111100001101010: color_data = 8'b11111111;
		20'b00010111100001101011: color_data = 8'b11111111;
		20'b00010111100001101100: color_data = 8'b11111111;
		20'b00010111100001101101: color_data = 8'b11111111;
		20'b00010111100001101110: color_data = 8'b11111111;
		20'b00010111100001101111: color_data = 8'b11111111;
		20'b00010111100001110000: color_data = 8'b11111111;
		20'b00010111100001110001: color_data = 8'b11111111;
		20'b00010111100001110010: color_data = 8'b10010010;
		20'b00010111100010000101: color_data = 8'b11011011;
		20'b00010111100010000110: color_data = 8'b11111111;
		20'b00010111100010000111: color_data = 8'b11111111;
		20'b00010111100010001000: color_data = 8'b11111111;
		20'b00010111100010001001: color_data = 8'b11111111;
		20'b00010111100010001010: color_data = 8'b11111111;
		20'b00010111100010001011: color_data = 8'b11111111;
		20'b00010111100010001100: color_data = 8'b11111111;
		20'b00010111100010001101: color_data = 8'b11111111;
		20'b00010111100010001110: color_data = 8'b11111111;
		20'b00010111100010011000: color_data = 8'b11011011;
		20'b00010111100010011001: color_data = 8'b11111111;
		20'b00010111100010011010: color_data = 8'b11111111;
		20'b00010111100010011011: color_data = 8'b11111111;
		20'b00010111100010011100: color_data = 8'b11111111;
		20'b00010111100010011101: color_data = 8'b11111111;
		20'b00010111100010011110: color_data = 8'b11111111;
		20'b00010111100010011111: color_data = 8'b11111111;
		20'b00010111100010100000: color_data = 8'b11111111;
		20'b00010111100010100001: color_data = 8'b11011011;

		20'b00010111110000001001: color_data = 8'b11011011;
		20'b00010111110000001010: color_data = 8'b11111111;
		20'b00010111110000001011: color_data = 8'b11111111;
		20'b00010111110000001100: color_data = 8'b11111111;
		20'b00010111110000001101: color_data = 8'b11111111;
		20'b00010111110000001110: color_data = 8'b11111111;
		20'b00010111110000001111: color_data = 8'b11111111;
		20'b00010111110000010000: color_data = 8'b11111111;
		20'b00010111110000010001: color_data = 8'b11111111;
		20'b00010111110000010010: color_data = 8'b11111111;
		20'b00010111110000010011: color_data = 8'b11011011;
		20'b00010111110000010100: color_data = 8'b11011011;
		20'b00010111110000010101: color_data = 8'b11011011;
		20'b00010111110000010110: color_data = 8'b11011011;
		20'b00010111110000010111: color_data = 8'b11011011;
		20'b00010111110000011000: color_data = 8'b11011011;
		20'b00010111110000011001: color_data = 8'b11011011;
		20'b00010111110000011010: color_data = 8'b11011011;
		20'b00010111110000011011: color_data = 8'b11011011;
		20'b00010111110000011100: color_data = 8'b11011011;
		20'b00010111110000011101: color_data = 8'b11011011;
		20'b00010111110000011110: color_data = 8'b11011011;
		20'b00010111110000011111: color_data = 8'b11011011;
		20'b00010111110000100000: color_data = 8'b11011011;
		20'b00010111110000100001: color_data = 8'b11011011;
		20'b00010111110000100010: color_data = 8'b11011011;
		20'b00010111110000100011: color_data = 8'b11011011;
		20'b00010111110000100100: color_data = 8'b11011011;
		20'b00010111110000100101: color_data = 8'b11011011;
		20'b00010111110000100110: color_data = 8'b11111111;
		20'b00010111110000100111: color_data = 8'b11111111;
		20'b00010111110000101000: color_data = 8'b11111111;
		20'b00010111110000101001: color_data = 8'b11111111;
		20'b00010111110000101010: color_data = 8'b11111111;
		20'b00010111110000101011: color_data = 8'b11111111;
		20'b00010111110000101100: color_data = 8'b11111111;
		20'b00010111110000101101: color_data = 8'b11111111;
		20'b00010111110000101110: color_data = 8'b11111111;
		20'b00010111110000101111: color_data = 8'b11011011;
		20'b00010111110000111001: color_data = 8'b11111111;
		20'b00010111110000111010: color_data = 8'b11111111;
		20'b00010111110000111011: color_data = 8'b11111111;
		20'b00010111110000111100: color_data = 8'b11111111;
		20'b00010111110000111101: color_data = 8'b11111111;
		20'b00010111110000111110: color_data = 8'b11111111;
		20'b00010111110000111111: color_data = 8'b11111111;
		20'b00010111110001000000: color_data = 8'b11111111;
		20'b00010111110001000001: color_data = 8'b11111111;
		20'b00010111110001000010: color_data = 8'b11011011;
		20'b00010111110001010101: color_data = 8'b10010010;
		20'b00010111110001010110: color_data = 8'b11111111;
		20'b00010111110001010111: color_data = 8'b11111111;
		20'b00010111110001011000: color_data = 8'b11111111;
		20'b00010111110001011001: color_data = 8'b11111111;
		20'b00010111110001011010: color_data = 8'b11111111;
		20'b00010111110001011011: color_data = 8'b11111111;
		20'b00010111110001011100: color_data = 8'b11111111;
		20'b00010111110001011101: color_data = 8'b11111111;
		20'b00010111110001011110: color_data = 8'b11111111;
		20'b00010111110001011111: color_data = 8'b10010010;
		20'b00010111110001101000: color_data = 8'b10010010;
		20'b00010111110001101001: color_data = 8'b11111111;
		20'b00010111110001101010: color_data = 8'b11111111;
		20'b00010111110001101011: color_data = 8'b11111111;
		20'b00010111110001101100: color_data = 8'b11111111;
		20'b00010111110001101101: color_data = 8'b11111111;
		20'b00010111110001101110: color_data = 8'b11111111;
		20'b00010111110001101111: color_data = 8'b11111111;
		20'b00010111110001110000: color_data = 8'b11111111;
		20'b00010111110001110001: color_data = 8'b11111111;
		20'b00010111110001110010: color_data = 8'b10010010;
		20'b00010111110010000101: color_data = 8'b11011011;
		20'b00010111110010000110: color_data = 8'b11111111;
		20'b00010111110010000111: color_data = 8'b11111111;
		20'b00010111110010001000: color_data = 8'b11111111;
		20'b00010111110010001001: color_data = 8'b11111111;
		20'b00010111110010001010: color_data = 8'b11111111;
		20'b00010111110010001011: color_data = 8'b11111111;
		20'b00010111110010001100: color_data = 8'b11111111;
		20'b00010111110010001101: color_data = 8'b11111111;
		20'b00010111110010001110: color_data = 8'b11111111;
		20'b00010111110010011000: color_data = 8'b11011011;
		20'b00010111110010011001: color_data = 8'b11111111;
		20'b00010111110010011010: color_data = 8'b11111111;
		20'b00010111110010011011: color_data = 8'b11111111;
		20'b00010111110010011100: color_data = 8'b11111111;
		20'b00010111110010011101: color_data = 8'b11111111;
		20'b00010111110010011110: color_data = 8'b11111111;
		20'b00010111110010011111: color_data = 8'b11111111;
		20'b00010111110010100000: color_data = 8'b11111111;
		20'b00010111110010100001: color_data = 8'b11011011;
		20'b00010111110010101011: color_data = 8'b10010010;
		20'b00010111110010101100: color_data = 8'b11011011;
		20'b00010111110010101101: color_data = 8'b11011011;
		20'b00010111110010101110: color_data = 8'b11011011;
		20'b00010111110010101111: color_data = 8'b11011011;
		20'b00010111110010110000: color_data = 8'b11011011;
		20'b00010111110010110001: color_data = 8'b11011011;
		20'b00010111110010110010: color_data = 8'b11011011;
		20'b00010111110010110011: color_data = 8'b11011011;
		20'b00010111110010110100: color_data = 8'b11011011;
		20'b00010111110010110101: color_data = 8'b11011011;
		20'b00010111110010110110: color_data = 8'b11011011;
		20'b00010111110010110111: color_data = 8'b11011011;
		20'b00010111110010111000: color_data = 8'b11011011;
		20'b00010111110010111001: color_data = 8'b11011011;
		20'b00010111110010111010: color_data = 8'b11011011;
		20'b00010111110010111011: color_data = 8'b11011011;
		20'b00010111110010111100: color_data = 8'b11011011;
		20'b00010111110010111101: color_data = 8'b11011011;
		20'b00010111110010111110: color_data = 8'b10010010;

		20'b00011000000000001001: color_data = 8'b11011011;
		20'b00011000000000001010: color_data = 8'b11111111;
		20'b00011000000000001011: color_data = 8'b11111111;
		20'b00011000000000001100: color_data = 8'b11111111;
		20'b00011000000000001101: color_data = 8'b11111111;
		20'b00011000000000001110: color_data = 8'b11111111;
		20'b00011000000000001111: color_data = 8'b11111111;
		20'b00011000000000010000: color_data = 8'b11111111;
		20'b00011000000000010001: color_data = 8'b11111111;
		20'b00011000000000010010: color_data = 8'b11111111;
		20'b00011000000000010011: color_data = 8'b11111111;
		20'b00011000000000010100: color_data = 8'b11111111;
		20'b00011000000000010101: color_data = 8'b11111111;
		20'b00011000000000010110: color_data = 8'b11111111;
		20'b00011000000000010111: color_data = 8'b11111111;
		20'b00011000000000011000: color_data = 8'b11111111;
		20'b00011000000000011001: color_data = 8'b11111111;
		20'b00011000000000011010: color_data = 8'b11111111;
		20'b00011000000000011011: color_data = 8'b11111111;
		20'b00011000000000011100: color_data = 8'b11111111;
		20'b00011000000000011101: color_data = 8'b11111111;
		20'b00011000000000011110: color_data = 8'b11111111;
		20'b00011000000000011111: color_data = 8'b11111111;
		20'b00011000000000100000: color_data = 8'b11111111;
		20'b00011000000000100001: color_data = 8'b11111111;
		20'b00011000000000100010: color_data = 8'b11111111;
		20'b00011000000000100011: color_data = 8'b11111111;
		20'b00011000000000100100: color_data = 8'b11111111;
		20'b00011000000000100101: color_data = 8'b11111111;
		20'b00011000000000100110: color_data = 8'b11111111;
		20'b00011000000000100111: color_data = 8'b11111111;
		20'b00011000000000101000: color_data = 8'b11111111;
		20'b00011000000000101001: color_data = 8'b11111111;
		20'b00011000000000101010: color_data = 8'b11111111;
		20'b00011000000000101011: color_data = 8'b11111111;
		20'b00011000000000101100: color_data = 8'b11111111;
		20'b00011000000000101101: color_data = 8'b11111111;
		20'b00011000000000101110: color_data = 8'b11111111;
		20'b00011000000000101111: color_data = 8'b11011011;
		20'b00011000000000111001: color_data = 8'b11111111;
		20'b00011000000000111010: color_data = 8'b11111111;
		20'b00011000000000111011: color_data = 8'b11111111;
		20'b00011000000000111100: color_data = 8'b11111111;
		20'b00011000000000111101: color_data = 8'b11111111;
		20'b00011000000000111110: color_data = 8'b11111111;
		20'b00011000000000111111: color_data = 8'b11111111;
		20'b00011000000001000000: color_data = 8'b11111111;
		20'b00011000000001000001: color_data = 8'b11111111;
		20'b00011000000001000010: color_data = 8'b11011011;
		20'b00011000000001010101: color_data = 8'b10010010;
		20'b00011000000001010110: color_data = 8'b11111111;
		20'b00011000000001010111: color_data = 8'b11111111;
		20'b00011000000001011000: color_data = 8'b11111111;
		20'b00011000000001011001: color_data = 8'b11111111;
		20'b00011000000001011010: color_data = 8'b11111111;
		20'b00011000000001011011: color_data = 8'b11111111;
		20'b00011000000001011100: color_data = 8'b11111111;
		20'b00011000000001011101: color_data = 8'b11111111;
		20'b00011000000001011110: color_data = 8'b11111111;
		20'b00011000000001011111: color_data = 8'b10010010;
		20'b00011000000001101000: color_data = 8'b10010010;
		20'b00011000000001101001: color_data = 8'b11111111;
		20'b00011000000001101010: color_data = 8'b11111111;
		20'b00011000000001101011: color_data = 8'b11111111;
		20'b00011000000001101100: color_data = 8'b11111111;
		20'b00011000000001101101: color_data = 8'b11111111;
		20'b00011000000001101110: color_data = 8'b11111111;
		20'b00011000000001101111: color_data = 8'b11111111;
		20'b00011000000001110000: color_data = 8'b11111111;
		20'b00011000000001110001: color_data = 8'b11111111;
		20'b00011000000001110010: color_data = 8'b10010010;
		20'b00011000000010000101: color_data = 8'b11011011;
		20'b00011000000010000110: color_data = 8'b11111111;
		20'b00011000000010000111: color_data = 8'b11111111;
		20'b00011000000010001000: color_data = 8'b11111111;
		20'b00011000000010001001: color_data = 8'b11111111;
		20'b00011000000010001010: color_data = 8'b11111111;
		20'b00011000000010001011: color_data = 8'b11111111;
		20'b00011000000010001100: color_data = 8'b11111111;
		20'b00011000000010001101: color_data = 8'b11111111;
		20'b00011000000010001110: color_data = 8'b11111111;
		20'b00011000000010011000: color_data = 8'b11011011;
		20'b00011000000010011001: color_data = 8'b11111111;
		20'b00011000000010011010: color_data = 8'b11111111;
		20'b00011000000010011011: color_data = 8'b11111111;
		20'b00011000000010011100: color_data = 8'b11111111;
		20'b00011000000010011101: color_data = 8'b11111111;
		20'b00011000000010011110: color_data = 8'b11111111;
		20'b00011000000010011111: color_data = 8'b11111111;
		20'b00011000000010100000: color_data = 8'b11111111;
		20'b00011000000010100001: color_data = 8'b11011011;
		20'b00011000000010101011: color_data = 8'b11011011;
		20'b00011000000010101100: color_data = 8'b11111111;
		20'b00011000000010101101: color_data = 8'b11111111;
		20'b00011000000010101110: color_data = 8'b11111111;
		20'b00011000000010101111: color_data = 8'b11111111;
		20'b00011000000010110000: color_data = 8'b11111111;
		20'b00011000000010110001: color_data = 8'b11111111;
		20'b00011000000010110010: color_data = 8'b11111111;
		20'b00011000000010110011: color_data = 8'b11111111;
		20'b00011000000010110100: color_data = 8'b11111111;
		20'b00011000000010110101: color_data = 8'b11111111;
		20'b00011000000010110110: color_data = 8'b11111111;
		20'b00011000000010110111: color_data = 8'b11111111;
		20'b00011000000010111000: color_data = 8'b11111111;
		20'b00011000000010111001: color_data = 8'b11111111;
		20'b00011000000010111010: color_data = 8'b11111111;
		20'b00011000000010111011: color_data = 8'b11111111;
		20'b00011000000010111100: color_data = 8'b11111111;
		20'b00011000000010111101: color_data = 8'b11111111;
		20'b00011000000010111110: color_data = 8'b11011011;

		20'b00011000010000001001: color_data = 8'b11011011;
		20'b00011000010000001010: color_data = 8'b11111111;
		20'b00011000010000001011: color_data = 8'b11111111;
		20'b00011000010000001100: color_data = 8'b11111111;
		20'b00011000010000001101: color_data = 8'b11111111;
		20'b00011000010000001110: color_data = 8'b11111111;
		20'b00011000010000001111: color_data = 8'b11111111;
		20'b00011000010000010000: color_data = 8'b11111111;
		20'b00011000010000010001: color_data = 8'b11111111;
		20'b00011000010000010010: color_data = 8'b11111111;
		20'b00011000010000010011: color_data = 8'b11111111;
		20'b00011000010000010100: color_data = 8'b11111111;
		20'b00011000010000010101: color_data = 8'b11111111;
		20'b00011000010000010110: color_data = 8'b11111111;
		20'b00011000010000010111: color_data = 8'b11111111;
		20'b00011000010000011000: color_data = 8'b11111111;
		20'b00011000010000011001: color_data = 8'b11111111;
		20'b00011000010000011010: color_data = 8'b11111111;
		20'b00011000010000011011: color_data = 8'b11111111;
		20'b00011000010000011100: color_data = 8'b11111111;
		20'b00011000010000011101: color_data = 8'b11111111;
		20'b00011000010000011110: color_data = 8'b11111111;
		20'b00011000010000011111: color_data = 8'b11111111;
		20'b00011000010000100000: color_data = 8'b11111111;
		20'b00011000010000100001: color_data = 8'b11111111;
		20'b00011000010000100010: color_data = 8'b11111111;
		20'b00011000010000100011: color_data = 8'b11111111;
		20'b00011000010000100100: color_data = 8'b11111111;
		20'b00011000010000100101: color_data = 8'b11111111;
		20'b00011000010000100110: color_data = 8'b11111111;
		20'b00011000010000100111: color_data = 8'b11111111;
		20'b00011000010000101000: color_data = 8'b11111111;
		20'b00011000010000101001: color_data = 8'b11111111;
		20'b00011000010000101010: color_data = 8'b11111111;
		20'b00011000010000101011: color_data = 8'b11111111;
		20'b00011000010000101100: color_data = 8'b11111111;
		20'b00011000010000101101: color_data = 8'b11111111;
		20'b00011000010000101110: color_data = 8'b11111111;
		20'b00011000010000101111: color_data = 8'b11011011;
		20'b00011000010000111001: color_data = 8'b11111111;
		20'b00011000010000111010: color_data = 8'b11111111;
		20'b00011000010000111011: color_data = 8'b11111111;
		20'b00011000010000111100: color_data = 8'b11111111;
		20'b00011000010000111101: color_data = 8'b11111111;
		20'b00011000010000111110: color_data = 8'b11111111;
		20'b00011000010000111111: color_data = 8'b11111111;
		20'b00011000010001000000: color_data = 8'b11111111;
		20'b00011000010001000001: color_data = 8'b11111111;
		20'b00011000010001000010: color_data = 8'b11011011;
		20'b00011000010001010101: color_data = 8'b10010010;
		20'b00011000010001010110: color_data = 8'b11111111;
		20'b00011000010001010111: color_data = 8'b11111111;
		20'b00011000010001011000: color_data = 8'b11111111;
		20'b00011000010001011001: color_data = 8'b11111111;
		20'b00011000010001011010: color_data = 8'b11111111;
		20'b00011000010001011011: color_data = 8'b11111111;
		20'b00011000010001011100: color_data = 8'b11111111;
		20'b00011000010001011101: color_data = 8'b11111111;
		20'b00011000010001011110: color_data = 8'b11111111;
		20'b00011000010001011111: color_data = 8'b10010010;
		20'b00011000010001101000: color_data = 8'b10010010;
		20'b00011000010001101001: color_data = 8'b11111111;
		20'b00011000010001101010: color_data = 8'b11111111;
		20'b00011000010001101011: color_data = 8'b11111111;
		20'b00011000010001101100: color_data = 8'b11111111;
		20'b00011000010001101101: color_data = 8'b11111111;
		20'b00011000010001101110: color_data = 8'b11111111;
		20'b00011000010001101111: color_data = 8'b11111111;
		20'b00011000010001110000: color_data = 8'b11111111;
		20'b00011000010001110001: color_data = 8'b11111111;
		20'b00011000010001110010: color_data = 8'b10010010;
		20'b00011000010010000101: color_data = 8'b11011011;
		20'b00011000010010000110: color_data = 8'b11111111;
		20'b00011000010010000111: color_data = 8'b11111111;
		20'b00011000010010001000: color_data = 8'b11111111;
		20'b00011000010010001001: color_data = 8'b11111111;
		20'b00011000010010001010: color_data = 8'b11111111;
		20'b00011000010010001011: color_data = 8'b11111111;
		20'b00011000010010001100: color_data = 8'b11111111;
		20'b00011000010010001101: color_data = 8'b11111111;
		20'b00011000010010001110: color_data = 8'b11111111;
		20'b00011000010010011000: color_data = 8'b11011011;
		20'b00011000010010011001: color_data = 8'b11111111;
		20'b00011000010010011010: color_data = 8'b11111111;
		20'b00011000010010011011: color_data = 8'b11111111;
		20'b00011000010010011100: color_data = 8'b11111111;
		20'b00011000010010011101: color_data = 8'b11111111;
		20'b00011000010010011110: color_data = 8'b11111111;
		20'b00011000010010011111: color_data = 8'b11111111;
		20'b00011000010010100000: color_data = 8'b11111111;
		20'b00011000010010100001: color_data = 8'b11011011;
		20'b00011000010010101011: color_data = 8'b11011011;
		20'b00011000010010101100: color_data = 8'b11111111;
		20'b00011000010010101101: color_data = 8'b11111111;
		20'b00011000010010101110: color_data = 8'b11111111;
		20'b00011000010010101111: color_data = 8'b11111111;
		20'b00011000010010110000: color_data = 8'b11111111;
		20'b00011000010010110001: color_data = 8'b11111111;
		20'b00011000010010110010: color_data = 8'b11111111;
		20'b00011000010010110011: color_data = 8'b11111111;
		20'b00011000010010110100: color_data = 8'b11111111;
		20'b00011000010010110101: color_data = 8'b11111111;
		20'b00011000010010110110: color_data = 8'b11111111;
		20'b00011000010010110111: color_data = 8'b11111111;
		20'b00011000010010111000: color_data = 8'b11111111;
		20'b00011000010010111001: color_data = 8'b11111111;
		20'b00011000010010111010: color_data = 8'b11111111;
		20'b00011000010010111011: color_data = 8'b11111111;
		20'b00011000010010111100: color_data = 8'b11111111;
		20'b00011000010010111101: color_data = 8'b11111111;
		20'b00011000010010111110: color_data = 8'b11011011;

		20'b00011000100000001001: color_data = 8'b11011011;
		20'b00011000100000001010: color_data = 8'b11111111;
		20'b00011000100000001011: color_data = 8'b11111111;
		20'b00011000100000001100: color_data = 8'b11111111;
		20'b00011000100000001101: color_data = 8'b11111111;
		20'b00011000100000001110: color_data = 8'b11111111;
		20'b00011000100000001111: color_data = 8'b11111111;
		20'b00011000100000010000: color_data = 8'b11111111;
		20'b00011000100000010001: color_data = 8'b11111111;
		20'b00011000100000010010: color_data = 8'b11111111;
		20'b00011000100000010011: color_data = 8'b11111111;
		20'b00011000100000010100: color_data = 8'b11111111;
		20'b00011000100000010101: color_data = 8'b11111111;
		20'b00011000100000010110: color_data = 8'b11111111;
		20'b00011000100000010111: color_data = 8'b11111111;
		20'b00011000100000011000: color_data = 8'b11111111;
		20'b00011000100000011001: color_data = 8'b11111111;
		20'b00011000100000011010: color_data = 8'b11111111;
		20'b00011000100000011011: color_data = 8'b11111111;
		20'b00011000100000011100: color_data = 8'b11111111;
		20'b00011000100000011101: color_data = 8'b11111111;
		20'b00011000100000011110: color_data = 8'b11111111;
		20'b00011000100000011111: color_data = 8'b11111111;
		20'b00011000100000100000: color_data = 8'b11111111;
		20'b00011000100000100001: color_data = 8'b11111111;
		20'b00011000100000100010: color_data = 8'b11111111;
		20'b00011000100000100011: color_data = 8'b11111111;
		20'b00011000100000100100: color_data = 8'b11111111;
		20'b00011000100000100101: color_data = 8'b11111111;
		20'b00011000100000100110: color_data = 8'b11111111;
		20'b00011000100000100111: color_data = 8'b11111111;
		20'b00011000100000101000: color_data = 8'b11111111;
		20'b00011000100000101001: color_data = 8'b11111111;
		20'b00011000100000101010: color_data = 8'b11111111;
		20'b00011000100000101011: color_data = 8'b11111111;
		20'b00011000100000101100: color_data = 8'b11111111;
		20'b00011000100000101101: color_data = 8'b11111111;
		20'b00011000100000101110: color_data = 8'b11111111;
		20'b00011000100000101111: color_data = 8'b11011011;
		20'b00011000100000111001: color_data = 8'b11111111;
		20'b00011000100000111010: color_data = 8'b11111111;
		20'b00011000100000111011: color_data = 8'b11111111;
		20'b00011000100000111100: color_data = 8'b11111111;
		20'b00011000100000111101: color_data = 8'b11111111;
		20'b00011000100000111110: color_data = 8'b11111111;
		20'b00011000100000111111: color_data = 8'b11111111;
		20'b00011000100001000000: color_data = 8'b11111111;
		20'b00011000100001000001: color_data = 8'b11111111;
		20'b00011000100001000010: color_data = 8'b11011011;
		20'b00011000100001010101: color_data = 8'b10010010;
		20'b00011000100001010110: color_data = 8'b11111111;
		20'b00011000100001010111: color_data = 8'b11111111;
		20'b00011000100001011000: color_data = 8'b11111111;
		20'b00011000100001011001: color_data = 8'b11111111;
		20'b00011000100001011010: color_data = 8'b11111111;
		20'b00011000100001011011: color_data = 8'b11111111;
		20'b00011000100001011100: color_data = 8'b11111111;
		20'b00011000100001011101: color_data = 8'b11111111;
		20'b00011000100001011110: color_data = 8'b11111111;
		20'b00011000100001011111: color_data = 8'b10010010;
		20'b00011000100001101000: color_data = 8'b10010010;
		20'b00011000100001101001: color_data = 8'b11111111;
		20'b00011000100001101010: color_data = 8'b11111111;
		20'b00011000100001101011: color_data = 8'b11111111;
		20'b00011000100001101100: color_data = 8'b11111111;
		20'b00011000100001101101: color_data = 8'b11111111;
		20'b00011000100001101110: color_data = 8'b11111111;
		20'b00011000100001101111: color_data = 8'b11111111;
		20'b00011000100001110000: color_data = 8'b11111111;
		20'b00011000100001110001: color_data = 8'b11111111;
		20'b00011000100001110010: color_data = 8'b10010010;
		20'b00011000100010000101: color_data = 8'b11011011;
		20'b00011000100010000110: color_data = 8'b11111111;
		20'b00011000100010000111: color_data = 8'b11111111;
		20'b00011000100010001000: color_data = 8'b11111111;
		20'b00011000100010001001: color_data = 8'b11111111;
		20'b00011000100010001010: color_data = 8'b11111111;
		20'b00011000100010001011: color_data = 8'b11111111;
		20'b00011000100010001100: color_data = 8'b11111111;
		20'b00011000100010001101: color_data = 8'b11111111;
		20'b00011000100010001110: color_data = 8'b11111111;
		20'b00011000100010011000: color_data = 8'b11011011;
		20'b00011000100010011001: color_data = 8'b11111111;
		20'b00011000100010011010: color_data = 8'b11111111;
		20'b00011000100010011011: color_data = 8'b11111111;
		20'b00011000100010011100: color_data = 8'b11111111;
		20'b00011000100010011101: color_data = 8'b11111111;
		20'b00011000100010011110: color_data = 8'b11111111;
		20'b00011000100010011111: color_data = 8'b11111111;
		20'b00011000100010100000: color_data = 8'b11111111;
		20'b00011000100010100001: color_data = 8'b11011011;
		20'b00011000100010101011: color_data = 8'b11011011;
		20'b00011000100010101100: color_data = 8'b11111111;
		20'b00011000100010101101: color_data = 8'b11111111;
		20'b00011000100010101110: color_data = 8'b11111111;
		20'b00011000100010101111: color_data = 8'b11111111;
		20'b00011000100010110000: color_data = 8'b11111111;
		20'b00011000100010110001: color_data = 8'b11111111;
		20'b00011000100010110010: color_data = 8'b11111111;
		20'b00011000100010110011: color_data = 8'b11111111;
		20'b00011000100010110100: color_data = 8'b11111111;
		20'b00011000100010110101: color_data = 8'b11111111;
		20'b00011000100010110110: color_data = 8'b11111111;
		20'b00011000100010110111: color_data = 8'b11111111;
		20'b00011000100010111000: color_data = 8'b11111111;
		20'b00011000100010111001: color_data = 8'b11111111;
		20'b00011000100010111010: color_data = 8'b11111111;
		20'b00011000100010111011: color_data = 8'b11111111;
		20'b00011000100010111100: color_data = 8'b11111111;
		20'b00011000100010111101: color_data = 8'b11111111;
		20'b00011000100010111110: color_data = 8'b11011011;

		20'b00011000110000001001: color_data = 8'b11011011;
		20'b00011000110000001010: color_data = 8'b11111111;
		20'b00011000110000001011: color_data = 8'b11111111;
		20'b00011000110000001100: color_data = 8'b11111111;
		20'b00011000110000001101: color_data = 8'b11111111;
		20'b00011000110000001110: color_data = 8'b11111111;
		20'b00011000110000001111: color_data = 8'b11111111;
		20'b00011000110000010000: color_data = 8'b11111111;
		20'b00011000110000010001: color_data = 8'b11111111;
		20'b00011000110000010010: color_data = 8'b11111111;
		20'b00011000110000010011: color_data = 8'b11111111;
		20'b00011000110000010100: color_data = 8'b11111111;
		20'b00011000110000010101: color_data = 8'b11111111;
		20'b00011000110000010110: color_data = 8'b11111111;
		20'b00011000110000010111: color_data = 8'b11111111;
		20'b00011000110000011000: color_data = 8'b11111111;
		20'b00011000110000011001: color_data = 8'b11111111;
		20'b00011000110000011010: color_data = 8'b11111111;
		20'b00011000110000011011: color_data = 8'b11111111;
		20'b00011000110000011100: color_data = 8'b11111111;
		20'b00011000110000011101: color_data = 8'b11111111;
		20'b00011000110000011110: color_data = 8'b11111111;
		20'b00011000110000011111: color_data = 8'b11111111;
		20'b00011000110000100000: color_data = 8'b11111111;
		20'b00011000110000100001: color_data = 8'b11111111;
		20'b00011000110000100010: color_data = 8'b11111111;
		20'b00011000110000100011: color_data = 8'b11111111;
		20'b00011000110000100100: color_data = 8'b11111111;
		20'b00011000110000100101: color_data = 8'b11111111;
		20'b00011000110000100110: color_data = 8'b11111111;
		20'b00011000110000100111: color_data = 8'b11111111;
		20'b00011000110000101000: color_data = 8'b11111111;
		20'b00011000110000101001: color_data = 8'b11111111;
		20'b00011000110000101010: color_data = 8'b11111111;
		20'b00011000110000101011: color_data = 8'b11111111;
		20'b00011000110000101100: color_data = 8'b11111111;
		20'b00011000110000101101: color_data = 8'b11111111;
		20'b00011000110000101110: color_data = 8'b11111111;
		20'b00011000110000101111: color_data = 8'b11011011;
		20'b00011000110000111001: color_data = 8'b11111111;
		20'b00011000110000111010: color_data = 8'b11111111;
		20'b00011000110000111011: color_data = 8'b11111111;
		20'b00011000110000111100: color_data = 8'b11111111;
		20'b00011000110000111101: color_data = 8'b11111111;
		20'b00011000110000111110: color_data = 8'b11111111;
		20'b00011000110000111111: color_data = 8'b11111111;
		20'b00011000110001000000: color_data = 8'b11111111;
		20'b00011000110001000001: color_data = 8'b11111111;
		20'b00011000110001000010: color_data = 8'b11011011;
		20'b00011000110001010101: color_data = 8'b10010010;
		20'b00011000110001010110: color_data = 8'b11111111;
		20'b00011000110001010111: color_data = 8'b11111111;
		20'b00011000110001011000: color_data = 8'b11111111;
		20'b00011000110001011001: color_data = 8'b11111111;
		20'b00011000110001011010: color_data = 8'b11111111;
		20'b00011000110001011011: color_data = 8'b11111111;
		20'b00011000110001011100: color_data = 8'b11111111;
		20'b00011000110001011101: color_data = 8'b11111111;
		20'b00011000110001011110: color_data = 8'b11111111;
		20'b00011000110001011111: color_data = 8'b10010010;
		20'b00011000110001101000: color_data = 8'b10010010;
		20'b00011000110001101001: color_data = 8'b11111111;
		20'b00011000110001101010: color_data = 8'b11111111;
		20'b00011000110001101011: color_data = 8'b11111111;
		20'b00011000110001101100: color_data = 8'b11111111;
		20'b00011000110001101101: color_data = 8'b11111111;
		20'b00011000110001101110: color_data = 8'b11111111;
		20'b00011000110001101111: color_data = 8'b11111111;
		20'b00011000110001110000: color_data = 8'b11111111;
		20'b00011000110001110001: color_data = 8'b11111111;
		20'b00011000110001110010: color_data = 8'b10010010;
		20'b00011000110010000101: color_data = 8'b11011011;
		20'b00011000110010000110: color_data = 8'b11111111;
		20'b00011000110010000111: color_data = 8'b11111111;
		20'b00011000110010001000: color_data = 8'b11111111;
		20'b00011000110010001001: color_data = 8'b11111111;
		20'b00011000110010001010: color_data = 8'b11111111;
		20'b00011000110010001011: color_data = 8'b11111111;
		20'b00011000110010001100: color_data = 8'b11111111;
		20'b00011000110010001101: color_data = 8'b11111111;
		20'b00011000110010001110: color_data = 8'b11111111;
		20'b00011000110010011000: color_data = 8'b11011011;
		20'b00011000110010011001: color_data = 8'b11111111;
		20'b00011000110010011010: color_data = 8'b11111111;
		20'b00011000110010011011: color_data = 8'b11111111;
		20'b00011000110010011100: color_data = 8'b11111111;
		20'b00011000110010011101: color_data = 8'b11111111;
		20'b00011000110010011110: color_data = 8'b11111111;
		20'b00011000110010011111: color_data = 8'b11111111;
		20'b00011000110010100000: color_data = 8'b11111111;
		20'b00011000110010100001: color_data = 8'b11011011;
		20'b00011000110010101011: color_data = 8'b11011011;
		20'b00011000110010101100: color_data = 8'b11111111;
		20'b00011000110010101101: color_data = 8'b11111111;
		20'b00011000110010101110: color_data = 8'b11111111;
		20'b00011000110010101111: color_data = 8'b11111111;
		20'b00011000110010110000: color_data = 8'b11111111;
		20'b00011000110010110001: color_data = 8'b11111111;
		20'b00011000110010110010: color_data = 8'b11111111;
		20'b00011000110010110011: color_data = 8'b11111111;
		20'b00011000110010110100: color_data = 8'b11111111;
		20'b00011000110010110101: color_data = 8'b11111111;
		20'b00011000110010110110: color_data = 8'b11111111;
		20'b00011000110010110111: color_data = 8'b11111111;
		20'b00011000110010111000: color_data = 8'b11111111;
		20'b00011000110010111001: color_data = 8'b11111111;
		20'b00011000110010111010: color_data = 8'b11111111;
		20'b00011000110010111011: color_data = 8'b11111111;
		20'b00011000110010111100: color_data = 8'b11111111;
		20'b00011000110010111101: color_data = 8'b11111111;
		20'b00011000110010111110: color_data = 8'b11011011;

		20'b00011001000000001001: color_data = 8'b11011011;
		20'b00011001000000001010: color_data = 8'b11111111;
		20'b00011001000000001011: color_data = 8'b11111111;
		20'b00011001000000001100: color_data = 8'b11111111;
		20'b00011001000000001101: color_data = 8'b11111111;
		20'b00011001000000001110: color_data = 8'b11111111;
		20'b00011001000000001111: color_data = 8'b11111111;
		20'b00011001000000010000: color_data = 8'b11111111;
		20'b00011001000000010001: color_data = 8'b11111111;
		20'b00011001000000010010: color_data = 8'b11111111;
		20'b00011001000000010011: color_data = 8'b11111111;
		20'b00011001000000010100: color_data = 8'b11111111;
		20'b00011001000000010101: color_data = 8'b11111111;
		20'b00011001000000010110: color_data = 8'b11111111;
		20'b00011001000000010111: color_data = 8'b11111111;
		20'b00011001000000011000: color_data = 8'b11111111;
		20'b00011001000000011001: color_data = 8'b11111111;
		20'b00011001000000011010: color_data = 8'b11111111;
		20'b00011001000000011011: color_data = 8'b11111111;
		20'b00011001000000011100: color_data = 8'b11111111;
		20'b00011001000000011101: color_data = 8'b11111111;
		20'b00011001000000011110: color_data = 8'b11111111;
		20'b00011001000000011111: color_data = 8'b11111111;
		20'b00011001000000100000: color_data = 8'b11111111;
		20'b00011001000000100001: color_data = 8'b11111111;
		20'b00011001000000100010: color_data = 8'b11111111;
		20'b00011001000000100011: color_data = 8'b11111111;
		20'b00011001000000100100: color_data = 8'b11111111;
		20'b00011001000000100101: color_data = 8'b11111111;
		20'b00011001000000100110: color_data = 8'b11111111;
		20'b00011001000000100111: color_data = 8'b11111111;
		20'b00011001000000101000: color_data = 8'b11111111;
		20'b00011001000000101001: color_data = 8'b11111111;
		20'b00011001000000101010: color_data = 8'b11111111;
		20'b00011001000000101011: color_data = 8'b11111111;
		20'b00011001000000101100: color_data = 8'b11111111;
		20'b00011001000000101101: color_data = 8'b11111111;
		20'b00011001000000101110: color_data = 8'b11111111;
		20'b00011001000000101111: color_data = 8'b11011011;
		20'b00011001000000111001: color_data = 8'b11111111;
		20'b00011001000000111010: color_data = 8'b11111111;
		20'b00011001000000111011: color_data = 8'b11111111;
		20'b00011001000000111100: color_data = 8'b11111111;
		20'b00011001000000111101: color_data = 8'b11111111;
		20'b00011001000000111110: color_data = 8'b11111111;
		20'b00011001000000111111: color_data = 8'b11111111;
		20'b00011001000001000000: color_data = 8'b11111111;
		20'b00011001000001000001: color_data = 8'b11111111;
		20'b00011001000001000010: color_data = 8'b11011011;
		20'b00011001000001010101: color_data = 8'b10010010;
		20'b00011001000001010110: color_data = 8'b11111111;
		20'b00011001000001010111: color_data = 8'b11111111;
		20'b00011001000001011000: color_data = 8'b11111111;
		20'b00011001000001011001: color_data = 8'b11111111;
		20'b00011001000001011010: color_data = 8'b11111111;
		20'b00011001000001011011: color_data = 8'b11111111;
		20'b00011001000001011100: color_data = 8'b11111111;
		20'b00011001000001011101: color_data = 8'b11111111;
		20'b00011001000001011110: color_data = 8'b11111111;
		20'b00011001000001011111: color_data = 8'b10010010;
		20'b00011001000001101000: color_data = 8'b10010010;
		20'b00011001000001101001: color_data = 8'b11111111;
		20'b00011001000001101010: color_data = 8'b11111111;
		20'b00011001000001101011: color_data = 8'b11111111;
		20'b00011001000001101100: color_data = 8'b11111111;
		20'b00011001000001101101: color_data = 8'b11111111;
		20'b00011001000001101110: color_data = 8'b11111111;
		20'b00011001000001101111: color_data = 8'b11111111;
		20'b00011001000001110000: color_data = 8'b11111111;
		20'b00011001000001110001: color_data = 8'b11111111;
		20'b00011001000001110010: color_data = 8'b10010010;
		20'b00011001000010000101: color_data = 8'b11011011;
		20'b00011001000010000110: color_data = 8'b11111111;
		20'b00011001000010000111: color_data = 8'b11111111;
		20'b00011001000010001000: color_data = 8'b11111111;
		20'b00011001000010001001: color_data = 8'b11111111;
		20'b00011001000010001010: color_data = 8'b11111111;
		20'b00011001000010001011: color_data = 8'b11111111;
		20'b00011001000010001100: color_data = 8'b11111111;
		20'b00011001000010001101: color_data = 8'b11111111;
		20'b00011001000010001110: color_data = 8'b11111111;
		20'b00011001000010011000: color_data = 8'b11011011;
		20'b00011001000010011001: color_data = 8'b11111111;
		20'b00011001000010011010: color_data = 8'b11111111;
		20'b00011001000010011011: color_data = 8'b11111111;
		20'b00011001000010011100: color_data = 8'b11111111;
		20'b00011001000010011101: color_data = 8'b11111111;
		20'b00011001000010011110: color_data = 8'b11111111;
		20'b00011001000010011111: color_data = 8'b11111111;
		20'b00011001000010100000: color_data = 8'b11111111;
		20'b00011001000010100001: color_data = 8'b11011011;
		20'b00011001000010101011: color_data = 8'b11011011;
		20'b00011001000010101100: color_data = 8'b11111111;
		20'b00011001000010101101: color_data = 8'b11111111;
		20'b00011001000010101110: color_data = 8'b11111111;
		20'b00011001000010101111: color_data = 8'b11111111;
		20'b00011001000010110000: color_data = 8'b11111111;
		20'b00011001000010110001: color_data = 8'b11111111;
		20'b00011001000010110010: color_data = 8'b11111111;
		20'b00011001000010110011: color_data = 8'b11111111;
		20'b00011001000010110100: color_data = 8'b11111111;
		20'b00011001000010110101: color_data = 8'b11111111;
		20'b00011001000010110110: color_data = 8'b11111111;
		20'b00011001000010110111: color_data = 8'b11111111;
		20'b00011001000010111000: color_data = 8'b11111111;
		20'b00011001000010111001: color_data = 8'b11111111;
		20'b00011001000010111010: color_data = 8'b11111111;
		20'b00011001000010111011: color_data = 8'b11111111;
		20'b00011001000010111100: color_data = 8'b11111111;
		20'b00011001000010111101: color_data = 8'b11111111;
		20'b00011001000010111110: color_data = 8'b11011011;

		20'b00011001010000001001: color_data = 8'b11011011;
		20'b00011001010000001010: color_data = 8'b11111111;
		20'b00011001010000001011: color_data = 8'b11111111;
		20'b00011001010000001100: color_data = 8'b11111111;
		20'b00011001010000001101: color_data = 8'b11111111;
		20'b00011001010000001110: color_data = 8'b11111111;
		20'b00011001010000001111: color_data = 8'b11111111;
		20'b00011001010000010000: color_data = 8'b11111111;
		20'b00011001010000010001: color_data = 8'b11111111;
		20'b00011001010000010010: color_data = 8'b11111111;
		20'b00011001010000010011: color_data = 8'b11111111;
		20'b00011001010000010100: color_data = 8'b11111111;
		20'b00011001010000010101: color_data = 8'b11111111;
		20'b00011001010000010110: color_data = 8'b11111111;
		20'b00011001010000010111: color_data = 8'b11111111;
		20'b00011001010000011000: color_data = 8'b11111111;
		20'b00011001010000011001: color_data = 8'b11111111;
		20'b00011001010000011010: color_data = 8'b11111111;
		20'b00011001010000011011: color_data = 8'b11111111;
		20'b00011001010000011100: color_data = 8'b11111111;
		20'b00011001010000011101: color_data = 8'b11111111;
		20'b00011001010000011110: color_data = 8'b11111111;
		20'b00011001010000011111: color_data = 8'b11111111;
		20'b00011001010000100000: color_data = 8'b11111111;
		20'b00011001010000100001: color_data = 8'b11111111;
		20'b00011001010000100010: color_data = 8'b11111111;
		20'b00011001010000100011: color_data = 8'b11111111;
		20'b00011001010000100100: color_data = 8'b11111111;
		20'b00011001010000100101: color_data = 8'b11111111;
		20'b00011001010000100110: color_data = 8'b11111111;
		20'b00011001010000100111: color_data = 8'b11111111;
		20'b00011001010000101000: color_data = 8'b11111111;
		20'b00011001010000101001: color_data = 8'b11111111;
		20'b00011001010000101010: color_data = 8'b11111111;
		20'b00011001010000101011: color_data = 8'b11111111;
		20'b00011001010000101100: color_data = 8'b11111111;
		20'b00011001010000101101: color_data = 8'b11111111;
		20'b00011001010000101110: color_data = 8'b11111111;
		20'b00011001010000101111: color_data = 8'b11011011;
		20'b00011001010000111001: color_data = 8'b11111111;
		20'b00011001010000111010: color_data = 8'b11111111;
		20'b00011001010000111011: color_data = 8'b11111111;
		20'b00011001010000111100: color_data = 8'b11111111;
		20'b00011001010000111101: color_data = 8'b11111111;
		20'b00011001010000111110: color_data = 8'b11111111;
		20'b00011001010000111111: color_data = 8'b11111111;
		20'b00011001010001000000: color_data = 8'b11111111;
		20'b00011001010001000001: color_data = 8'b11111111;
		20'b00011001010001000010: color_data = 8'b11011011;
		20'b00011001010001010101: color_data = 8'b10010010;
		20'b00011001010001010110: color_data = 8'b11111111;
		20'b00011001010001010111: color_data = 8'b11111111;
		20'b00011001010001011000: color_data = 8'b11111111;
		20'b00011001010001011001: color_data = 8'b11111111;
		20'b00011001010001011010: color_data = 8'b11111111;
		20'b00011001010001011011: color_data = 8'b11111111;
		20'b00011001010001011100: color_data = 8'b11111111;
		20'b00011001010001011101: color_data = 8'b11111111;
		20'b00011001010001011110: color_data = 8'b11111111;
		20'b00011001010001011111: color_data = 8'b10010010;
		20'b00011001010001101000: color_data = 8'b10010010;
		20'b00011001010001101001: color_data = 8'b11111111;
		20'b00011001010001101010: color_data = 8'b11111111;
		20'b00011001010001101011: color_data = 8'b11111111;
		20'b00011001010001101100: color_data = 8'b11111111;
		20'b00011001010001101101: color_data = 8'b11111111;
		20'b00011001010001101110: color_data = 8'b11111111;
		20'b00011001010001101111: color_data = 8'b11111111;
		20'b00011001010001110000: color_data = 8'b11111111;
		20'b00011001010001110001: color_data = 8'b11111111;
		20'b00011001010001110010: color_data = 8'b10010010;
		20'b00011001010010000101: color_data = 8'b11011011;
		20'b00011001010010000110: color_data = 8'b11111111;
		20'b00011001010010000111: color_data = 8'b11111111;
		20'b00011001010010001000: color_data = 8'b11111111;
		20'b00011001010010001001: color_data = 8'b11111111;
		20'b00011001010010001010: color_data = 8'b11111111;
		20'b00011001010010001011: color_data = 8'b11111111;
		20'b00011001010010001100: color_data = 8'b11111111;
		20'b00011001010010001101: color_data = 8'b11111111;
		20'b00011001010010001110: color_data = 8'b11111111;
		20'b00011001010010011000: color_data = 8'b11011011;
		20'b00011001010010011001: color_data = 8'b11111111;
		20'b00011001010010011010: color_data = 8'b11111111;
		20'b00011001010010011011: color_data = 8'b11111111;
		20'b00011001010010011100: color_data = 8'b11111111;
		20'b00011001010010011101: color_data = 8'b11111111;
		20'b00011001010010011110: color_data = 8'b11111111;
		20'b00011001010010011111: color_data = 8'b11111111;
		20'b00011001010010100000: color_data = 8'b11111111;
		20'b00011001010010100001: color_data = 8'b11011011;
		20'b00011001010010101011: color_data = 8'b11011011;
		20'b00011001010010101100: color_data = 8'b11111111;
		20'b00011001010010101101: color_data = 8'b11111111;
		20'b00011001010010101110: color_data = 8'b11111111;
		20'b00011001010010101111: color_data = 8'b11111111;
		20'b00011001010010110000: color_data = 8'b11111111;
		20'b00011001010010110001: color_data = 8'b11111111;
		20'b00011001010010110010: color_data = 8'b11111111;
		20'b00011001010010110011: color_data = 8'b11111111;
		20'b00011001010010110100: color_data = 8'b11111111;
		20'b00011001010010110101: color_data = 8'b11111111;
		20'b00011001010010110110: color_data = 8'b11111111;
		20'b00011001010010110111: color_data = 8'b11111111;
		20'b00011001010010111000: color_data = 8'b11111111;
		20'b00011001010010111001: color_data = 8'b11111111;
		20'b00011001010010111010: color_data = 8'b11111111;
		20'b00011001010010111011: color_data = 8'b11111111;
		20'b00011001010010111100: color_data = 8'b11111111;
		20'b00011001010010111101: color_data = 8'b11111111;
		20'b00011001010010111110: color_data = 8'b11011011;

		20'b00011001100000001001: color_data = 8'b11011011;
		20'b00011001100000001010: color_data = 8'b11111111;
		20'b00011001100000001011: color_data = 8'b11111111;
		20'b00011001100000001100: color_data = 8'b11111111;
		20'b00011001100000001101: color_data = 8'b11111111;
		20'b00011001100000001110: color_data = 8'b11111111;
		20'b00011001100000001111: color_data = 8'b11111111;
		20'b00011001100000010000: color_data = 8'b11111111;
		20'b00011001100000010001: color_data = 8'b11111111;
		20'b00011001100000010010: color_data = 8'b11111111;
		20'b00011001100000010011: color_data = 8'b11111111;
		20'b00011001100000010100: color_data = 8'b11111111;
		20'b00011001100000010101: color_data = 8'b11111111;
		20'b00011001100000010110: color_data = 8'b11111111;
		20'b00011001100000010111: color_data = 8'b11111111;
		20'b00011001100000011000: color_data = 8'b11111111;
		20'b00011001100000011001: color_data = 8'b11111111;
		20'b00011001100000011010: color_data = 8'b11111111;
		20'b00011001100000011011: color_data = 8'b11111111;
		20'b00011001100000011100: color_data = 8'b11111111;
		20'b00011001100000011101: color_data = 8'b11111111;
		20'b00011001100000011110: color_data = 8'b11111111;
		20'b00011001100000011111: color_data = 8'b11111111;
		20'b00011001100000100000: color_data = 8'b11111111;
		20'b00011001100000100001: color_data = 8'b11111111;
		20'b00011001100000100010: color_data = 8'b11111111;
		20'b00011001100000100011: color_data = 8'b11111111;
		20'b00011001100000100100: color_data = 8'b11111111;
		20'b00011001100000100101: color_data = 8'b11111111;
		20'b00011001100000100110: color_data = 8'b11111111;
		20'b00011001100000100111: color_data = 8'b11111111;
		20'b00011001100000101000: color_data = 8'b11111111;
		20'b00011001100000101001: color_data = 8'b11111111;
		20'b00011001100000101010: color_data = 8'b11111111;
		20'b00011001100000101011: color_data = 8'b11111111;
		20'b00011001100000101100: color_data = 8'b11111111;
		20'b00011001100000101101: color_data = 8'b11111111;
		20'b00011001100000101110: color_data = 8'b11111111;
		20'b00011001100000101111: color_data = 8'b11011011;
		20'b00011001100000111001: color_data = 8'b11111111;
		20'b00011001100000111010: color_data = 8'b11111111;
		20'b00011001100000111011: color_data = 8'b11111111;
		20'b00011001100000111100: color_data = 8'b11111111;
		20'b00011001100000111101: color_data = 8'b11111111;
		20'b00011001100000111110: color_data = 8'b11111111;
		20'b00011001100000111111: color_data = 8'b11111111;
		20'b00011001100001000000: color_data = 8'b11111111;
		20'b00011001100001000001: color_data = 8'b11111111;
		20'b00011001100001000010: color_data = 8'b11011011;
		20'b00011001100001010101: color_data = 8'b10010010;
		20'b00011001100001010110: color_data = 8'b11111111;
		20'b00011001100001010111: color_data = 8'b11111111;
		20'b00011001100001011000: color_data = 8'b11111111;
		20'b00011001100001011001: color_data = 8'b11111111;
		20'b00011001100001011010: color_data = 8'b11111111;
		20'b00011001100001011011: color_data = 8'b11111111;
		20'b00011001100001011100: color_data = 8'b11111111;
		20'b00011001100001011101: color_data = 8'b11111111;
		20'b00011001100001011110: color_data = 8'b11111111;
		20'b00011001100001011111: color_data = 8'b10010010;
		20'b00011001100001101000: color_data = 8'b10010010;
		20'b00011001100001101001: color_data = 8'b11111111;
		20'b00011001100001101010: color_data = 8'b11111111;
		20'b00011001100001101011: color_data = 8'b11111111;
		20'b00011001100001101100: color_data = 8'b11111111;
		20'b00011001100001101101: color_data = 8'b11111111;
		20'b00011001100001101110: color_data = 8'b11111111;
		20'b00011001100001101111: color_data = 8'b11111111;
		20'b00011001100001110000: color_data = 8'b11111111;
		20'b00011001100001110001: color_data = 8'b11111111;
		20'b00011001100001110010: color_data = 8'b10010010;
		20'b00011001100010000101: color_data = 8'b11011011;
		20'b00011001100010000110: color_data = 8'b11111111;
		20'b00011001100010000111: color_data = 8'b11111111;
		20'b00011001100010001000: color_data = 8'b11111111;
		20'b00011001100010001001: color_data = 8'b11111111;
		20'b00011001100010001010: color_data = 8'b11111111;
		20'b00011001100010001011: color_data = 8'b11111111;
		20'b00011001100010001100: color_data = 8'b11111111;
		20'b00011001100010001101: color_data = 8'b11111111;
		20'b00011001100010001110: color_data = 8'b11111111;
		20'b00011001100010011000: color_data = 8'b11011011;
		20'b00011001100010011001: color_data = 8'b11111111;
		20'b00011001100010011010: color_data = 8'b11111111;
		20'b00011001100010011011: color_data = 8'b11111111;
		20'b00011001100010011100: color_data = 8'b11111111;
		20'b00011001100010011101: color_data = 8'b11111111;
		20'b00011001100010011110: color_data = 8'b11111111;
		20'b00011001100010011111: color_data = 8'b11111111;
		20'b00011001100010100000: color_data = 8'b11111111;
		20'b00011001100010100001: color_data = 8'b11011011;
		20'b00011001100010101011: color_data = 8'b11011011;
		20'b00011001100010101100: color_data = 8'b11111111;
		20'b00011001100010101101: color_data = 8'b11111111;
		20'b00011001100010101110: color_data = 8'b11111111;
		20'b00011001100010101111: color_data = 8'b11111111;
		20'b00011001100010110000: color_data = 8'b11111111;
		20'b00011001100010110001: color_data = 8'b11111111;
		20'b00011001100010110010: color_data = 8'b11111111;
		20'b00011001100010110011: color_data = 8'b11111111;
		20'b00011001100010110100: color_data = 8'b11111111;
		20'b00011001100010110101: color_data = 8'b11111111;
		20'b00011001100010110110: color_data = 8'b11111111;
		20'b00011001100010110111: color_data = 8'b11111111;
		20'b00011001100010111000: color_data = 8'b11111111;
		20'b00011001100010111001: color_data = 8'b11111111;
		20'b00011001100010111010: color_data = 8'b11111111;
		20'b00011001100010111011: color_data = 8'b11111111;
		20'b00011001100010111100: color_data = 8'b11111111;
		20'b00011001100010111101: color_data = 8'b11111111;
		20'b00011001100010111110: color_data = 8'b11011011;

		20'b00011001110000001001: color_data = 8'b11011011;
		20'b00011001110000001010: color_data = 8'b11111111;
		20'b00011001110000001011: color_data = 8'b11111111;
		20'b00011001110000001100: color_data = 8'b11111111;
		20'b00011001110000001101: color_data = 8'b11111111;
		20'b00011001110000001110: color_data = 8'b11111111;
		20'b00011001110000001111: color_data = 8'b11111111;
		20'b00011001110000010000: color_data = 8'b11111111;
		20'b00011001110000010001: color_data = 8'b11111111;
		20'b00011001110000010010: color_data = 8'b11111111;
		20'b00011001110000010011: color_data = 8'b11111111;
		20'b00011001110000010100: color_data = 8'b11111111;
		20'b00011001110000010101: color_data = 8'b11111111;
		20'b00011001110000010110: color_data = 8'b11111111;
		20'b00011001110000010111: color_data = 8'b11111111;
		20'b00011001110000011000: color_data = 8'b11111111;
		20'b00011001110000011001: color_data = 8'b11111111;
		20'b00011001110000011010: color_data = 8'b11111111;
		20'b00011001110000011011: color_data = 8'b11111111;
		20'b00011001110000011100: color_data = 8'b11111111;
		20'b00011001110000011101: color_data = 8'b11111111;
		20'b00011001110000011110: color_data = 8'b11111111;
		20'b00011001110000011111: color_data = 8'b11111111;
		20'b00011001110000100000: color_data = 8'b11111111;
		20'b00011001110000100001: color_data = 8'b11111111;
		20'b00011001110000100010: color_data = 8'b11111111;
		20'b00011001110000100011: color_data = 8'b11111111;
		20'b00011001110000100100: color_data = 8'b11111111;
		20'b00011001110000100101: color_data = 8'b11111111;
		20'b00011001110000100110: color_data = 8'b11111111;
		20'b00011001110000100111: color_data = 8'b11111111;
		20'b00011001110000101000: color_data = 8'b11111111;
		20'b00011001110000101001: color_data = 8'b11111111;
		20'b00011001110000101010: color_data = 8'b11111111;
		20'b00011001110000101011: color_data = 8'b11111111;
		20'b00011001110000101100: color_data = 8'b11111111;
		20'b00011001110000101101: color_data = 8'b11111111;
		20'b00011001110000101110: color_data = 8'b11111111;
		20'b00011001110000101111: color_data = 8'b11011011;
		20'b00011001110000111001: color_data = 8'b11111111;
		20'b00011001110000111010: color_data = 8'b11111111;
		20'b00011001110000111011: color_data = 8'b11111111;
		20'b00011001110000111100: color_data = 8'b11111111;
		20'b00011001110000111101: color_data = 8'b11111111;
		20'b00011001110000111110: color_data = 8'b11111111;
		20'b00011001110000111111: color_data = 8'b11111111;
		20'b00011001110001000000: color_data = 8'b11111111;
		20'b00011001110001000001: color_data = 8'b11111111;
		20'b00011001110001000010: color_data = 8'b11011011;
		20'b00011001110001010101: color_data = 8'b10010010;
		20'b00011001110001010110: color_data = 8'b11111111;
		20'b00011001110001010111: color_data = 8'b11111111;
		20'b00011001110001011000: color_data = 8'b11111111;
		20'b00011001110001011001: color_data = 8'b11111111;
		20'b00011001110001011010: color_data = 8'b11111111;
		20'b00011001110001011011: color_data = 8'b11111111;
		20'b00011001110001011100: color_data = 8'b11111111;
		20'b00011001110001011101: color_data = 8'b11111111;
		20'b00011001110001011110: color_data = 8'b11111111;
		20'b00011001110001011111: color_data = 8'b10010010;
		20'b00011001110001101000: color_data = 8'b10010010;
		20'b00011001110001101001: color_data = 8'b11111111;
		20'b00011001110001101010: color_data = 8'b11111111;
		20'b00011001110001101011: color_data = 8'b11111111;
		20'b00011001110001101100: color_data = 8'b11111111;
		20'b00011001110001101101: color_data = 8'b11111111;
		20'b00011001110001101110: color_data = 8'b11111111;
		20'b00011001110001101111: color_data = 8'b11111111;
		20'b00011001110001110000: color_data = 8'b11111111;
		20'b00011001110001110001: color_data = 8'b11111111;
		20'b00011001110001110010: color_data = 8'b10010010;
		20'b00011001110010000101: color_data = 8'b11011011;
		20'b00011001110010000110: color_data = 8'b11111111;
		20'b00011001110010000111: color_data = 8'b11111111;
		20'b00011001110010001000: color_data = 8'b11111111;
		20'b00011001110010001001: color_data = 8'b11111111;
		20'b00011001110010001010: color_data = 8'b11111111;
		20'b00011001110010001011: color_data = 8'b11111111;
		20'b00011001110010001100: color_data = 8'b11111111;
		20'b00011001110010001101: color_data = 8'b11111111;
		20'b00011001110010001110: color_data = 8'b11111111;
		20'b00011001110010011000: color_data = 8'b11011011;
		20'b00011001110010011001: color_data = 8'b11111111;
		20'b00011001110010011010: color_data = 8'b11111111;
		20'b00011001110010011011: color_data = 8'b11111111;
		20'b00011001110010011100: color_data = 8'b11111111;
		20'b00011001110010011101: color_data = 8'b11111111;
		20'b00011001110010011110: color_data = 8'b11111111;
		20'b00011001110010011111: color_data = 8'b11111111;
		20'b00011001110010100000: color_data = 8'b11111111;
		20'b00011001110010100001: color_data = 8'b11011011;
		20'b00011001110010101011: color_data = 8'b11011011;
		20'b00011001110010101100: color_data = 8'b11111111;
		20'b00011001110010101101: color_data = 8'b11111111;
		20'b00011001110010101110: color_data = 8'b11111111;
		20'b00011001110010101111: color_data = 8'b11111111;
		20'b00011001110010110000: color_data = 8'b11111111;
		20'b00011001110010110001: color_data = 8'b11111111;
		20'b00011001110010110010: color_data = 8'b11111111;
		20'b00011001110010110011: color_data = 8'b11111111;
		20'b00011001110010110100: color_data = 8'b11111111;
		20'b00011001110010110101: color_data = 8'b11111111;
		20'b00011001110010110110: color_data = 8'b11111111;
		20'b00011001110010110111: color_data = 8'b11111111;
		20'b00011001110010111000: color_data = 8'b11111111;
		20'b00011001110010111001: color_data = 8'b11111111;
		20'b00011001110010111010: color_data = 8'b11111111;
		20'b00011001110010111011: color_data = 8'b11111111;
		20'b00011001110010111100: color_data = 8'b11111111;
		20'b00011001110010111101: color_data = 8'b11111111;
		20'b00011001110010111110: color_data = 8'b11011011;

		20'b00011010000000001001: color_data = 8'b11011011;
		20'b00011010000000001010: color_data = 8'b11111111;
		20'b00011010000000001011: color_data = 8'b11111111;
		20'b00011010000000001100: color_data = 8'b11111111;
		20'b00011010000000001101: color_data = 8'b11111111;
		20'b00011010000000001110: color_data = 8'b11111111;
		20'b00011010000000001111: color_data = 8'b11111111;
		20'b00011010000000010000: color_data = 8'b11111111;
		20'b00011010000000010001: color_data = 8'b11111111;
		20'b00011010000000010010: color_data = 8'b11111111;
		20'b00011010000000010011: color_data = 8'b11011011;
		20'b00011010000000010100: color_data = 8'b11011011;
		20'b00011010000000010101: color_data = 8'b11011011;
		20'b00011010000000010110: color_data = 8'b11011011;
		20'b00011010000000010111: color_data = 8'b11011011;
		20'b00011010000000011000: color_data = 8'b11011011;
		20'b00011010000000011001: color_data = 8'b11011011;
		20'b00011010000000011010: color_data = 8'b11011011;
		20'b00011010000000011011: color_data = 8'b11011011;
		20'b00011010000000011100: color_data = 8'b11011011;
		20'b00011010000000011101: color_data = 8'b11011011;
		20'b00011010000000011110: color_data = 8'b11011011;
		20'b00011010000000011111: color_data = 8'b11011011;
		20'b00011010000000100000: color_data = 8'b11011011;
		20'b00011010000000100001: color_data = 8'b11011011;
		20'b00011010000000100010: color_data = 8'b11011011;
		20'b00011010000000100011: color_data = 8'b11011011;
		20'b00011010000000100100: color_data = 8'b11011011;
		20'b00011010000000100101: color_data = 8'b11011011;
		20'b00011010000000100110: color_data = 8'b11011011;
		20'b00011010000000100111: color_data = 8'b11011011;
		20'b00011010000000101000: color_data = 8'b11011011;
		20'b00011010000000101001: color_data = 8'b11011011;
		20'b00011010000000101010: color_data = 8'b11011011;
		20'b00011010000000101011: color_data = 8'b11011011;
		20'b00011010000000101100: color_data = 8'b11011011;
		20'b00011010000000101101: color_data = 8'b11011011;
		20'b00011010000000101110: color_data = 8'b11011011;
		20'b00011010000000101111: color_data = 8'b11011011;
		20'b00011010000000111001: color_data = 8'b11111111;
		20'b00011010000000111010: color_data = 8'b11111111;
		20'b00011010000000111011: color_data = 8'b11111111;
		20'b00011010000000111100: color_data = 8'b11111111;
		20'b00011010000000111101: color_data = 8'b11111111;
		20'b00011010000000111110: color_data = 8'b11111111;
		20'b00011010000000111111: color_data = 8'b11111111;
		20'b00011010000001000000: color_data = 8'b11111111;
		20'b00011010000001000001: color_data = 8'b11111111;
		20'b00011010000001000010: color_data = 8'b11011011;
		20'b00011010000001010101: color_data = 8'b10010010;
		20'b00011010000001010110: color_data = 8'b11111111;
		20'b00011010000001010111: color_data = 8'b11111111;
		20'b00011010000001011000: color_data = 8'b11111111;
		20'b00011010000001011001: color_data = 8'b11111111;
		20'b00011010000001011010: color_data = 8'b11111111;
		20'b00011010000001011011: color_data = 8'b11111111;
		20'b00011010000001011100: color_data = 8'b11111111;
		20'b00011010000001011101: color_data = 8'b11111111;
		20'b00011010000001011110: color_data = 8'b11111111;
		20'b00011010000001011111: color_data = 8'b10010010;
		20'b00011010000001101000: color_data = 8'b10010010;
		20'b00011010000001101001: color_data = 8'b11111111;
		20'b00011010000001101010: color_data = 8'b11111111;
		20'b00011010000001101011: color_data = 8'b11111111;
		20'b00011010000001101100: color_data = 8'b11111111;
		20'b00011010000001101101: color_data = 8'b11111111;
		20'b00011010000001101110: color_data = 8'b11111111;
		20'b00011010000001101111: color_data = 8'b11111111;
		20'b00011010000001110000: color_data = 8'b11111111;
		20'b00011010000001110001: color_data = 8'b11111111;
		20'b00011010000001110010: color_data = 8'b10010010;
		20'b00011010000010000101: color_data = 8'b11011011;
		20'b00011010000010000110: color_data = 8'b11111111;
		20'b00011010000010000111: color_data = 8'b11111111;
		20'b00011010000010001000: color_data = 8'b11111111;
		20'b00011010000010001001: color_data = 8'b11111111;
		20'b00011010000010001010: color_data = 8'b11111111;
		20'b00011010000010001011: color_data = 8'b11111111;
		20'b00011010000010001100: color_data = 8'b11111111;
		20'b00011010000010001101: color_data = 8'b11111111;
		20'b00011010000010001110: color_data = 8'b11111111;
		20'b00011010000010011000: color_data = 8'b11011011;
		20'b00011010000010011001: color_data = 8'b11111111;
		20'b00011010000010011010: color_data = 8'b11111111;
		20'b00011010000010011011: color_data = 8'b11111111;
		20'b00011010000010011100: color_data = 8'b11111111;
		20'b00011010000010011101: color_data = 8'b11111111;
		20'b00011010000010011110: color_data = 8'b11111111;
		20'b00011010000010011111: color_data = 8'b11111111;
		20'b00011010000010100000: color_data = 8'b11111111;
		20'b00011010000010100001: color_data = 8'b11011011;
		20'b00011010000010101011: color_data = 8'b10010010;
		20'b00011010000010101100: color_data = 8'b11011011;
		20'b00011010000010101101: color_data = 8'b11011011;
		20'b00011010000010101110: color_data = 8'b11011011;
		20'b00011010000010101111: color_data = 8'b11011011;
		20'b00011010000010110000: color_data = 8'b11011011;
		20'b00011010000010110001: color_data = 8'b11011011;
		20'b00011010000010110010: color_data = 8'b11011011;
		20'b00011010000010110011: color_data = 8'b11011011;
		20'b00011010000010110100: color_data = 8'b11011011;
		20'b00011010000010110101: color_data = 8'b11111111;
		20'b00011010000010110110: color_data = 8'b11111111;
		20'b00011010000010110111: color_data = 8'b11111111;
		20'b00011010000010111000: color_data = 8'b11111111;
		20'b00011010000010111001: color_data = 8'b11111111;
		20'b00011010000010111010: color_data = 8'b11111111;
		20'b00011010000010111011: color_data = 8'b11111111;
		20'b00011010000010111100: color_data = 8'b11111111;
		20'b00011010000010111101: color_data = 8'b11111111;
		20'b00011010000010111110: color_data = 8'b11011011;

		20'b00011010010000001001: color_data = 8'b11011011;
		20'b00011010010000001010: color_data = 8'b11111111;
		20'b00011010010000001011: color_data = 8'b11111111;
		20'b00011010010000001100: color_data = 8'b11111111;
		20'b00011010010000001101: color_data = 8'b11111111;
		20'b00011010010000001110: color_data = 8'b11111111;
		20'b00011010010000001111: color_data = 8'b11111111;
		20'b00011010010000010000: color_data = 8'b11111111;
		20'b00011010010000010001: color_data = 8'b11111111;
		20'b00011010010000010010: color_data = 8'b11111111;
		20'b00011010010000010011: color_data = 8'b10010010;
		20'b00011010010000111001: color_data = 8'b11111111;
		20'b00011010010000111010: color_data = 8'b11111111;
		20'b00011010010000111011: color_data = 8'b11111111;
		20'b00011010010000111100: color_data = 8'b11111111;
		20'b00011010010000111101: color_data = 8'b11111111;
		20'b00011010010000111110: color_data = 8'b11111111;
		20'b00011010010000111111: color_data = 8'b11111111;
		20'b00011010010001000000: color_data = 8'b11111111;
		20'b00011010010001000001: color_data = 8'b11111111;
		20'b00011010010001000010: color_data = 8'b11011011;
		20'b00011010010001010101: color_data = 8'b10010010;
		20'b00011010010001010110: color_data = 8'b11111111;
		20'b00011010010001010111: color_data = 8'b11111111;
		20'b00011010010001011000: color_data = 8'b11111111;
		20'b00011010010001011001: color_data = 8'b11111111;
		20'b00011010010001011010: color_data = 8'b11111111;
		20'b00011010010001011011: color_data = 8'b11111111;
		20'b00011010010001011100: color_data = 8'b11111111;
		20'b00011010010001011101: color_data = 8'b11111111;
		20'b00011010010001011110: color_data = 8'b11111111;
		20'b00011010010001011111: color_data = 8'b10010010;
		20'b00011010010001101000: color_data = 8'b10010010;
		20'b00011010010001101001: color_data = 8'b11111111;
		20'b00011010010001101010: color_data = 8'b11111111;
		20'b00011010010001101011: color_data = 8'b11111111;
		20'b00011010010001101100: color_data = 8'b11111111;
		20'b00011010010001101101: color_data = 8'b11111111;
		20'b00011010010001101110: color_data = 8'b11111111;
		20'b00011010010001101111: color_data = 8'b11111111;
		20'b00011010010001110000: color_data = 8'b11111111;
		20'b00011010010001110001: color_data = 8'b11111111;
		20'b00011010010001110010: color_data = 8'b10010010;
		20'b00011010010010000101: color_data = 8'b11011011;
		20'b00011010010010000110: color_data = 8'b11111111;
		20'b00011010010010000111: color_data = 8'b11111111;
		20'b00011010010010001000: color_data = 8'b11111111;
		20'b00011010010010001001: color_data = 8'b11111111;
		20'b00011010010010001010: color_data = 8'b11111111;
		20'b00011010010010001011: color_data = 8'b11111111;
		20'b00011010010010001100: color_data = 8'b11111111;
		20'b00011010010010001101: color_data = 8'b11111111;
		20'b00011010010010001110: color_data = 8'b11111111;
		20'b00011010010010011000: color_data = 8'b11011011;
		20'b00011010010010011001: color_data = 8'b11111111;
		20'b00011010010010011010: color_data = 8'b11111111;
		20'b00011010010010011011: color_data = 8'b11111111;
		20'b00011010010010011100: color_data = 8'b11111111;
		20'b00011010010010011101: color_data = 8'b11111111;
		20'b00011010010010011110: color_data = 8'b11111111;
		20'b00011010010010011111: color_data = 8'b11111111;
		20'b00011010010010100000: color_data = 8'b11111111;
		20'b00011010010010100001: color_data = 8'b11011011;
		20'b00011010010010110100: color_data = 8'b10010010;
		20'b00011010010010110101: color_data = 8'b11111111;
		20'b00011010010010110110: color_data = 8'b11111111;
		20'b00011010010010110111: color_data = 8'b11111111;
		20'b00011010010010111000: color_data = 8'b11111111;
		20'b00011010010010111001: color_data = 8'b11111111;
		20'b00011010010010111010: color_data = 8'b11111111;
		20'b00011010010010111011: color_data = 8'b11111111;
		20'b00011010010010111100: color_data = 8'b11111111;
		20'b00011010010010111101: color_data = 8'b11111111;
		20'b00011010010010111110: color_data = 8'b11011011;

		20'b00011010100000001001: color_data = 8'b11011011;
		20'b00011010100000001010: color_data = 8'b11111111;
		20'b00011010100000001011: color_data = 8'b11111111;
		20'b00011010100000001100: color_data = 8'b11111111;
		20'b00011010100000001101: color_data = 8'b11111111;
		20'b00011010100000001110: color_data = 8'b11111111;
		20'b00011010100000001111: color_data = 8'b11111111;
		20'b00011010100000010000: color_data = 8'b11111111;
		20'b00011010100000010001: color_data = 8'b11111111;
		20'b00011010100000010010: color_data = 8'b11111111;
		20'b00011010100000010011: color_data = 8'b10010010;
		20'b00011010100000111001: color_data = 8'b11111111;
		20'b00011010100000111010: color_data = 8'b11111111;
		20'b00011010100000111011: color_data = 8'b11111111;
		20'b00011010100000111100: color_data = 8'b11111111;
		20'b00011010100000111101: color_data = 8'b11111111;
		20'b00011010100000111110: color_data = 8'b11111111;
		20'b00011010100000111111: color_data = 8'b11111111;
		20'b00011010100001000000: color_data = 8'b11111111;
		20'b00011010100001000001: color_data = 8'b11111111;
		20'b00011010100001000010: color_data = 8'b11011011;
		20'b00011010100001010101: color_data = 8'b10010010;
		20'b00011010100001010110: color_data = 8'b11111111;
		20'b00011010100001010111: color_data = 8'b11111111;
		20'b00011010100001011000: color_data = 8'b11111111;
		20'b00011010100001011001: color_data = 8'b11111111;
		20'b00011010100001011010: color_data = 8'b11111111;
		20'b00011010100001011011: color_data = 8'b11111111;
		20'b00011010100001011100: color_data = 8'b11111111;
		20'b00011010100001011101: color_data = 8'b11111111;
		20'b00011010100001011110: color_data = 8'b11111111;
		20'b00011010100001011111: color_data = 8'b10010010;
		20'b00011010100001101000: color_data = 8'b10010010;
		20'b00011010100001101001: color_data = 8'b11111111;
		20'b00011010100001101010: color_data = 8'b11111111;
		20'b00011010100001101011: color_data = 8'b11111111;
		20'b00011010100001101100: color_data = 8'b11111111;
		20'b00011010100001101101: color_data = 8'b11111111;
		20'b00011010100001101110: color_data = 8'b11111111;
		20'b00011010100001101111: color_data = 8'b11111111;
		20'b00011010100001110000: color_data = 8'b11111111;
		20'b00011010100001110001: color_data = 8'b11111111;
		20'b00011010100001110010: color_data = 8'b10010010;
		20'b00011010100010000101: color_data = 8'b11011011;
		20'b00011010100010000110: color_data = 8'b11111111;
		20'b00011010100010000111: color_data = 8'b11111111;
		20'b00011010100010001000: color_data = 8'b11111111;
		20'b00011010100010001001: color_data = 8'b11111111;
		20'b00011010100010001010: color_data = 8'b11111111;
		20'b00011010100010001011: color_data = 8'b11111111;
		20'b00011010100010001100: color_data = 8'b11111111;
		20'b00011010100010001101: color_data = 8'b11111111;
		20'b00011010100010001110: color_data = 8'b11111111;
		20'b00011010100010011000: color_data = 8'b11011011;
		20'b00011010100010011001: color_data = 8'b11111111;
		20'b00011010100010011010: color_data = 8'b11111111;
		20'b00011010100010011011: color_data = 8'b11111111;
		20'b00011010100010011100: color_data = 8'b11111111;
		20'b00011010100010011101: color_data = 8'b11111111;
		20'b00011010100010011110: color_data = 8'b11111111;
		20'b00011010100010011111: color_data = 8'b11111111;
		20'b00011010100010100000: color_data = 8'b11111111;
		20'b00011010100010100001: color_data = 8'b11011011;
		20'b00011010100010110100: color_data = 8'b10010010;
		20'b00011010100010110101: color_data = 8'b11111111;
		20'b00011010100010110110: color_data = 8'b11111111;
		20'b00011010100010110111: color_data = 8'b11111111;
		20'b00011010100010111000: color_data = 8'b11111111;
		20'b00011010100010111001: color_data = 8'b11111111;
		20'b00011010100010111010: color_data = 8'b11111111;
		20'b00011010100010111011: color_data = 8'b11111111;
		20'b00011010100010111100: color_data = 8'b11111111;
		20'b00011010100010111101: color_data = 8'b11111111;
		20'b00011010100010111110: color_data = 8'b11011011;

		20'b00011010110000001001: color_data = 8'b11011011;
		20'b00011010110000001010: color_data = 8'b11111111;
		20'b00011010110000001011: color_data = 8'b11111111;
		20'b00011010110000001100: color_data = 8'b11111111;
		20'b00011010110000001101: color_data = 8'b11111111;
		20'b00011010110000001110: color_data = 8'b11111111;
		20'b00011010110000001111: color_data = 8'b11111111;
		20'b00011010110000010000: color_data = 8'b11111111;
		20'b00011010110000010001: color_data = 8'b11111111;
		20'b00011010110000010010: color_data = 8'b11111111;
		20'b00011010110000010011: color_data = 8'b10010010;
		20'b00011010110000111001: color_data = 8'b11111111;
		20'b00011010110000111010: color_data = 8'b11111111;
		20'b00011010110000111011: color_data = 8'b11111111;
		20'b00011010110000111100: color_data = 8'b11111111;
		20'b00011010110000111101: color_data = 8'b11111111;
		20'b00011010110000111110: color_data = 8'b11111111;
		20'b00011010110000111111: color_data = 8'b11111111;
		20'b00011010110001000000: color_data = 8'b11111111;
		20'b00011010110001000001: color_data = 8'b11111111;
		20'b00011010110001000010: color_data = 8'b11011011;
		20'b00011010110001010101: color_data = 8'b10010010;
		20'b00011010110001010110: color_data = 8'b11111111;
		20'b00011010110001010111: color_data = 8'b11111111;
		20'b00011010110001011000: color_data = 8'b11111111;
		20'b00011010110001011001: color_data = 8'b11111111;
		20'b00011010110001011010: color_data = 8'b11111111;
		20'b00011010110001011011: color_data = 8'b11111111;
		20'b00011010110001011100: color_data = 8'b11111111;
		20'b00011010110001011101: color_data = 8'b11111111;
		20'b00011010110001011110: color_data = 8'b11111111;
		20'b00011010110001011111: color_data = 8'b10010010;
		20'b00011010110001101000: color_data = 8'b10010010;
		20'b00011010110001101001: color_data = 8'b11111111;
		20'b00011010110001101010: color_data = 8'b11111111;
		20'b00011010110001101011: color_data = 8'b11111111;
		20'b00011010110001101100: color_data = 8'b11111111;
		20'b00011010110001101101: color_data = 8'b11111111;
		20'b00011010110001101110: color_data = 8'b11111111;
		20'b00011010110001101111: color_data = 8'b11111111;
		20'b00011010110001110000: color_data = 8'b11111111;
		20'b00011010110001110001: color_data = 8'b11111111;
		20'b00011010110001110010: color_data = 8'b10010010;
		20'b00011010110010000101: color_data = 8'b11011011;
		20'b00011010110010000110: color_data = 8'b11111111;
		20'b00011010110010000111: color_data = 8'b11111111;
		20'b00011010110010001000: color_data = 8'b11111111;
		20'b00011010110010001001: color_data = 8'b11111111;
		20'b00011010110010001010: color_data = 8'b11111111;
		20'b00011010110010001011: color_data = 8'b11111111;
		20'b00011010110010001100: color_data = 8'b11111111;
		20'b00011010110010001101: color_data = 8'b11111111;
		20'b00011010110010001110: color_data = 8'b11111111;
		20'b00011010110010011000: color_data = 8'b11011011;
		20'b00011010110010011001: color_data = 8'b11111111;
		20'b00011010110010011010: color_data = 8'b11111111;
		20'b00011010110010011011: color_data = 8'b11111111;
		20'b00011010110010011100: color_data = 8'b11111111;
		20'b00011010110010011101: color_data = 8'b11111111;
		20'b00011010110010011110: color_data = 8'b11111111;
		20'b00011010110010011111: color_data = 8'b11111111;
		20'b00011010110010100000: color_data = 8'b11111111;
		20'b00011010110010100001: color_data = 8'b11011011;
		20'b00011010110010110100: color_data = 8'b10010010;
		20'b00011010110010110101: color_data = 8'b11111111;
		20'b00011010110010110110: color_data = 8'b11111111;
		20'b00011010110010110111: color_data = 8'b11111111;
		20'b00011010110010111000: color_data = 8'b11111111;
		20'b00011010110010111001: color_data = 8'b11111111;
		20'b00011010110010111010: color_data = 8'b11111111;
		20'b00011010110010111011: color_data = 8'b11111111;
		20'b00011010110010111100: color_data = 8'b11111111;
		20'b00011010110010111101: color_data = 8'b11111111;
		20'b00011010110010111110: color_data = 8'b11011011;

		20'b00011011000000001001: color_data = 8'b11011011;
		20'b00011011000000001010: color_data = 8'b11111111;
		20'b00011011000000001011: color_data = 8'b11111111;
		20'b00011011000000001100: color_data = 8'b11111111;
		20'b00011011000000001101: color_data = 8'b11111111;
		20'b00011011000000001110: color_data = 8'b11111111;
		20'b00011011000000001111: color_data = 8'b11111111;
		20'b00011011000000010000: color_data = 8'b11111111;
		20'b00011011000000010001: color_data = 8'b11111111;
		20'b00011011000000010010: color_data = 8'b11111111;
		20'b00011011000000010011: color_data = 8'b10010010;
		20'b00011011000000111001: color_data = 8'b11111111;
		20'b00011011000000111010: color_data = 8'b11111111;
		20'b00011011000000111011: color_data = 8'b11111111;
		20'b00011011000000111100: color_data = 8'b11111111;
		20'b00011011000000111101: color_data = 8'b11111111;
		20'b00011011000000111110: color_data = 8'b11111111;
		20'b00011011000000111111: color_data = 8'b11111111;
		20'b00011011000001000000: color_data = 8'b11111111;
		20'b00011011000001000001: color_data = 8'b11111111;
		20'b00011011000001000010: color_data = 8'b11011011;
		20'b00011011000001010101: color_data = 8'b10010010;
		20'b00011011000001010110: color_data = 8'b11111111;
		20'b00011011000001010111: color_data = 8'b11111111;
		20'b00011011000001011000: color_data = 8'b11111111;
		20'b00011011000001011001: color_data = 8'b11111111;
		20'b00011011000001011010: color_data = 8'b11111111;
		20'b00011011000001011011: color_data = 8'b11111111;
		20'b00011011000001011100: color_data = 8'b11111111;
		20'b00011011000001011101: color_data = 8'b11111111;
		20'b00011011000001011110: color_data = 8'b11111111;
		20'b00011011000001011111: color_data = 8'b10010010;
		20'b00011011000001101000: color_data = 8'b10010010;
		20'b00011011000001101001: color_data = 8'b11111111;
		20'b00011011000001101010: color_data = 8'b11111111;
		20'b00011011000001101011: color_data = 8'b11111111;
		20'b00011011000001101100: color_data = 8'b11111111;
		20'b00011011000001101101: color_data = 8'b11111111;
		20'b00011011000001101110: color_data = 8'b11111111;
		20'b00011011000001101111: color_data = 8'b11111111;
		20'b00011011000001110000: color_data = 8'b11111111;
		20'b00011011000001110001: color_data = 8'b11111111;
		20'b00011011000001110010: color_data = 8'b10010010;
		20'b00011011000010000101: color_data = 8'b11011011;
		20'b00011011000010000110: color_data = 8'b11111111;
		20'b00011011000010000111: color_data = 8'b11111111;
		20'b00011011000010001000: color_data = 8'b11111111;
		20'b00011011000010001001: color_data = 8'b11111111;
		20'b00011011000010001010: color_data = 8'b11111111;
		20'b00011011000010001011: color_data = 8'b11111111;
		20'b00011011000010001100: color_data = 8'b11111111;
		20'b00011011000010001101: color_data = 8'b11111111;
		20'b00011011000010001110: color_data = 8'b11111111;
		20'b00011011000010011000: color_data = 8'b11011011;
		20'b00011011000010011001: color_data = 8'b11111111;
		20'b00011011000010011010: color_data = 8'b11111111;
		20'b00011011000010011011: color_data = 8'b11111111;
		20'b00011011000010011100: color_data = 8'b11111111;
		20'b00011011000010011101: color_data = 8'b11111111;
		20'b00011011000010011110: color_data = 8'b11111111;
		20'b00011011000010011111: color_data = 8'b11111111;
		20'b00011011000010100000: color_data = 8'b11111111;
		20'b00011011000010100001: color_data = 8'b11011011;
		20'b00011011000010110100: color_data = 8'b10010010;
		20'b00011011000010110101: color_data = 8'b11111111;
		20'b00011011000010110110: color_data = 8'b11111111;
		20'b00011011000010110111: color_data = 8'b11111111;
		20'b00011011000010111000: color_data = 8'b11111111;
		20'b00011011000010111001: color_data = 8'b11111111;
		20'b00011011000010111010: color_data = 8'b11111111;
		20'b00011011000010111011: color_data = 8'b11111111;
		20'b00011011000010111100: color_data = 8'b11111111;
		20'b00011011000010111101: color_data = 8'b11111111;
		20'b00011011000010111110: color_data = 8'b11011011;

		20'b00011011010000001001: color_data = 8'b11011011;
		20'b00011011010000001010: color_data = 8'b11111111;
		20'b00011011010000001011: color_data = 8'b11111111;
		20'b00011011010000001100: color_data = 8'b11111111;
		20'b00011011010000001101: color_data = 8'b11111111;
		20'b00011011010000001110: color_data = 8'b11111111;
		20'b00011011010000001111: color_data = 8'b11111111;
		20'b00011011010000010000: color_data = 8'b11111111;
		20'b00011011010000010001: color_data = 8'b11111111;
		20'b00011011010000010010: color_data = 8'b11111111;
		20'b00011011010000010011: color_data = 8'b10010010;
		20'b00011011010000111001: color_data = 8'b11111111;
		20'b00011011010000111010: color_data = 8'b11111111;
		20'b00011011010000111011: color_data = 8'b11111111;
		20'b00011011010000111100: color_data = 8'b11111111;
		20'b00011011010000111101: color_data = 8'b11111111;
		20'b00011011010000111110: color_data = 8'b11111111;
		20'b00011011010000111111: color_data = 8'b11111111;
		20'b00011011010001000000: color_data = 8'b11111111;
		20'b00011011010001000001: color_data = 8'b11111111;
		20'b00011011010001000010: color_data = 8'b11011011;
		20'b00011011010001010101: color_data = 8'b10010010;
		20'b00011011010001010110: color_data = 8'b11111111;
		20'b00011011010001010111: color_data = 8'b11111111;
		20'b00011011010001011000: color_data = 8'b11111111;
		20'b00011011010001011001: color_data = 8'b11111111;
		20'b00011011010001011010: color_data = 8'b11111111;
		20'b00011011010001011011: color_data = 8'b11111111;
		20'b00011011010001011100: color_data = 8'b11111111;
		20'b00011011010001011101: color_data = 8'b11111111;
		20'b00011011010001011110: color_data = 8'b11111111;
		20'b00011011010001011111: color_data = 8'b10010010;
		20'b00011011010001101000: color_data = 8'b10010010;
		20'b00011011010001101001: color_data = 8'b11111111;
		20'b00011011010001101010: color_data = 8'b11111111;
		20'b00011011010001101011: color_data = 8'b11111111;
		20'b00011011010001101100: color_data = 8'b11111111;
		20'b00011011010001101101: color_data = 8'b11111111;
		20'b00011011010001101110: color_data = 8'b11111111;
		20'b00011011010001101111: color_data = 8'b11111111;
		20'b00011011010001110000: color_data = 8'b11111111;
		20'b00011011010001110001: color_data = 8'b11111111;
		20'b00011011010001110010: color_data = 8'b10010010;
		20'b00011011010010000101: color_data = 8'b11011011;
		20'b00011011010010000110: color_data = 8'b11111111;
		20'b00011011010010000111: color_data = 8'b11111111;
		20'b00011011010010001000: color_data = 8'b11111111;
		20'b00011011010010001001: color_data = 8'b11111111;
		20'b00011011010010001010: color_data = 8'b11111111;
		20'b00011011010010001011: color_data = 8'b11111111;
		20'b00011011010010001100: color_data = 8'b11111111;
		20'b00011011010010001101: color_data = 8'b11111111;
		20'b00011011010010001110: color_data = 8'b11111111;
		20'b00011011010010011000: color_data = 8'b11011011;
		20'b00011011010010011001: color_data = 8'b11111111;
		20'b00011011010010011010: color_data = 8'b11111111;
		20'b00011011010010011011: color_data = 8'b11111111;
		20'b00011011010010011100: color_data = 8'b11111111;
		20'b00011011010010011101: color_data = 8'b11111111;
		20'b00011011010010011110: color_data = 8'b11111111;
		20'b00011011010010011111: color_data = 8'b11111111;
		20'b00011011010010100000: color_data = 8'b11111111;
		20'b00011011010010100001: color_data = 8'b11011011;
		20'b00011011010010110100: color_data = 8'b10010010;
		20'b00011011010010110101: color_data = 8'b11111111;
		20'b00011011010010110110: color_data = 8'b11111111;
		20'b00011011010010110111: color_data = 8'b11111111;
		20'b00011011010010111000: color_data = 8'b11111111;
		20'b00011011010010111001: color_data = 8'b11111111;
		20'b00011011010010111010: color_data = 8'b11111111;
		20'b00011011010010111011: color_data = 8'b11111111;
		20'b00011011010010111100: color_data = 8'b11111111;
		20'b00011011010010111101: color_data = 8'b11111111;
		20'b00011011010010111110: color_data = 8'b11011011;

		20'b00011011100000001001: color_data = 8'b11011011;
		20'b00011011100000001010: color_data = 8'b11111111;
		20'b00011011100000001011: color_data = 8'b11111111;
		20'b00011011100000001100: color_data = 8'b11111111;
		20'b00011011100000001101: color_data = 8'b11111111;
		20'b00011011100000001110: color_data = 8'b11111111;
		20'b00011011100000001111: color_data = 8'b11111111;
		20'b00011011100000010000: color_data = 8'b11111111;
		20'b00011011100000010001: color_data = 8'b11111111;
		20'b00011011100000010010: color_data = 8'b11111111;
		20'b00011011100000010011: color_data = 8'b10010010;
		20'b00011011100000111001: color_data = 8'b11111111;
		20'b00011011100000111010: color_data = 8'b11111111;
		20'b00011011100000111011: color_data = 8'b11111111;
		20'b00011011100000111100: color_data = 8'b11111111;
		20'b00011011100000111101: color_data = 8'b11111111;
		20'b00011011100000111110: color_data = 8'b11111111;
		20'b00011011100000111111: color_data = 8'b11111111;
		20'b00011011100001000000: color_data = 8'b11111111;
		20'b00011011100001000001: color_data = 8'b11111111;
		20'b00011011100001000010: color_data = 8'b11011011;
		20'b00011011100001010101: color_data = 8'b10010010;
		20'b00011011100001010110: color_data = 8'b11111111;
		20'b00011011100001010111: color_data = 8'b11111111;
		20'b00011011100001011000: color_data = 8'b11111111;
		20'b00011011100001011001: color_data = 8'b11111111;
		20'b00011011100001011010: color_data = 8'b11111111;
		20'b00011011100001011011: color_data = 8'b11111111;
		20'b00011011100001011100: color_data = 8'b11111111;
		20'b00011011100001011101: color_data = 8'b11111111;
		20'b00011011100001011110: color_data = 8'b11111111;
		20'b00011011100001011111: color_data = 8'b10010010;
		20'b00011011100001101000: color_data = 8'b10010010;
		20'b00011011100001101001: color_data = 8'b11111111;
		20'b00011011100001101010: color_data = 8'b11111111;
		20'b00011011100001101011: color_data = 8'b11111111;
		20'b00011011100001101100: color_data = 8'b11111111;
		20'b00011011100001101101: color_data = 8'b11111111;
		20'b00011011100001101110: color_data = 8'b11111111;
		20'b00011011100001101111: color_data = 8'b11111111;
		20'b00011011100001110000: color_data = 8'b11111111;
		20'b00011011100001110001: color_data = 8'b11111111;
		20'b00011011100001110010: color_data = 8'b10010010;
		20'b00011011100010000101: color_data = 8'b11011011;
		20'b00011011100010000110: color_data = 8'b11111111;
		20'b00011011100010000111: color_data = 8'b11111111;
		20'b00011011100010001000: color_data = 8'b11111111;
		20'b00011011100010001001: color_data = 8'b11111111;
		20'b00011011100010001010: color_data = 8'b11111111;
		20'b00011011100010001011: color_data = 8'b11111111;
		20'b00011011100010001100: color_data = 8'b11111111;
		20'b00011011100010001101: color_data = 8'b11111111;
		20'b00011011100010001110: color_data = 8'b11111111;
		20'b00011011100010011000: color_data = 8'b11011011;
		20'b00011011100010011001: color_data = 8'b11111111;
		20'b00011011100010011010: color_data = 8'b11111111;
		20'b00011011100010011011: color_data = 8'b11111111;
		20'b00011011100010011100: color_data = 8'b11111111;
		20'b00011011100010011101: color_data = 8'b11111111;
		20'b00011011100010011110: color_data = 8'b11111111;
		20'b00011011100010011111: color_data = 8'b11111111;
		20'b00011011100010100000: color_data = 8'b11111111;
		20'b00011011100010100001: color_data = 8'b11011011;
		20'b00011011100010110100: color_data = 8'b10010010;
		20'b00011011100010110101: color_data = 8'b11111111;
		20'b00011011100010110110: color_data = 8'b11111111;
		20'b00011011100010110111: color_data = 8'b11111111;
		20'b00011011100010111000: color_data = 8'b11111111;
		20'b00011011100010111001: color_data = 8'b11111111;
		20'b00011011100010111010: color_data = 8'b11111111;
		20'b00011011100010111011: color_data = 8'b11111111;
		20'b00011011100010111100: color_data = 8'b11111111;
		20'b00011011100010111101: color_data = 8'b11111111;
		20'b00011011100010111110: color_data = 8'b11011011;

		20'b00011011110000001001: color_data = 8'b11011011;
		20'b00011011110000001010: color_data = 8'b11111111;
		20'b00011011110000001011: color_data = 8'b11111111;
		20'b00011011110000001100: color_data = 8'b11111111;
		20'b00011011110000001101: color_data = 8'b11111111;
		20'b00011011110000001110: color_data = 8'b11111111;
		20'b00011011110000001111: color_data = 8'b11111111;
		20'b00011011110000010000: color_data = 8'b11111111;
		20'b00011011110000010001: color_data = 8'b11111111;
		20'b00011011110000010010: color_data = 8'b11111111;
		20'b00011011110000010011: color_data = 8'b10010010;
		20'b00011011110000111001: color_data = 8'b11111111;
		20'b00011011110000111010: color_data = 8'b11111111;
		20'b00011011110000111011: color_data = 8'b11111111;
		20'b00011011110000111100: color_data = 8'b11111111;
		20'b00011011110000111101: color_data = 8'b11111111;
		20'b00011011110000111110: color_data = 8'b11111111;
		20'b00011011110000111111: color_data = 8'b11111111;
		20'b00011011110001000000: color_data = 8'b11111111;
		20'b00011011110001000001: color_data = 8'b11111111;
		20'b00011011110001000010: color_data = 8'b11011011;
		20'b00011011110001010101: color_data = 8'b10010010;
		20'b00011011110001010110: color_data = 8'b11111111;
		20'b00011011110001010111: color_data = 8'b11111111;
		20'b00011011110001011000: color_data = 8'b11111111;
		20'b00011011110001011001: color_data = 8'b11111111;
		20'b00011011110001011010: color_data = 8'b11111111;
		20'b00011011110001011011: color_data = 8'b11111111;
		20'b00011011110001011100: color_data = 8'b11111111;
		20'b00011011110001011101: color_data = 8'b11111111;
		20'b00011011110001011110: color_data = 8'b11111111;
		20'b00011011110001011111: color_data = 8'b10010010;
		20'b00011011110001101000: color_data = 8'b10010010;
		20'b00011011110001101001: color_data = 8'b11111111;
		20'b00011011110001101010: color_data = 8'b11111111;
		20'b00011011110001101011: color_data = 8'b11111111;
		20'b00011011110001101100: color_data = 8'b11111111;
		20'b00011011110001101101: color_data = 8'b11111111;
		20'b00011011110001101110: color_data = 8'b11111111;
		20'b00011011110001101111: color_data = 8'b11111111;
		20'b00011011110001110000: color_data = 8'b11111111;
		20'b00011011110001110001: color_data = 8'b11111111;
		20'b00011011110001110010: color_data = 8'b10010010;
		20'b00011011110010000101: color_data = 8'b11011011;
		20'b00011011110010000110: color_data = 8'b11111111;
		20'b00011011110010000111: color_data = 8'b11111111;
		20'b00011011110010001000: color_data = 8'b11111111;
		20'b00011011110010001001: color_data = 8'b11111111;
		20'b00011011110010001010: color_data = 8'b11111111;
		20'b00011011110010001011: color_data = 8'b11111111;
		20'b00011011110010001100: color_data = 8'b11111111;
		20'b00011011110010001101: color_data = 8'b11111111;
		20'b00011011110010001110: color_data = 8'b11111111;
		20'b00011011110010011000: color_data = 8'b11011011;
		20'b00011011110010011001: color_data = 8'b11111111;
		20'b00011011110010011010: color_data = 8'b11111111;
		20'b00011011110010011011: color_data = 8'b11111111;
		20'b00011011110010011100: color_data = 8'b11111111;
		20'b00011011110010011101: color_data = 8'b11111111;
		20'b00011011110010011110: color_data = 8'b11111111;
		20'b00011011110010011111: color_data = 8'b11111111;
		20'b00011011110010100000: color_data = 8'b11111111;
		20'b00011011110010100001: color_data = 8'b11011011;
		20'b00011011110010110100: color_data = 8'b10010010;
		20'b00011011110010110101: color_data = 8'b11111111;
		20'b00011011110010110110: color_data = 8'b11111111;
		20'b00011011110010110111: color_data = 8'b11111111;
		20'b00011011110010111000: color_data = 8'b11111111;
		20'b00011011110010111001: color_data = 8'b11111111;
		20'b00011011110010111010: color_data = 8'b11111111;
		20'b00011011110010111011: color_data = 8'b11111111;
		20'b00011011110010111100: color_data = 8'b11111111;
		20'b00011011110010111101: color_data = 8'b11111111;
		20'b00011011110010111110: color_data = 8'b11011011;

		20'b00011100000000001001: color_data = 8'b11011011;
		20'b00011100000000001010: color_data = 8'b11111111;
		20'b00011100000000001011: color_data = 8'b11111111;
		20'b00011100000000001100: color_data = 8'b11111111;
		20'b00011100000000001101: color_data = 8'b11111111;
		20'b00011100000000001110: color_data = 8'b11111111;
		20'b00011100000000001111: color_data = 8'b11111111;
		20'b00011100000000010000: color_data = 8'b11111111;
		20'b00011100000000010001: color_data = 8'b11111111;
		20'b00011100000000010010: color_data = 8'b11111111;
		20'b00011100000000010011: color_data = 8'b10010010;
		20'b00011100000000111001: color_data = 8'b11111111;
		20'b00011100000000111010: color_data = 8'b11111111;
		20'b00011100000000111011: color_data = 8'b11111111;
		20'b00011100000000111100: color_data = 8'b11111111;
		20'b00011100000000111101: color_data = 8'b11111111;
		20'b00011100000000111110: color_data = 8'b11111111;
		20'b00011100000000111111: color_data = 8'b11111111;
		20'b00011100000001000000: color_data = 8'b11111111;
		20'b00011100000001000001: color_data = 8'b11111111;
		20'b00011100000001000010: color_data = 8'b11011011;
		20'b00011100000001010101: color_data = 8'b10010010;
		20'b00011100000001010110: color_data = 8'b11111111;
		20'b00011100000001010111: color_data = 8'b11111111;
		20'b00011100000001011000: color_data = 8'b11111111;
		20'b00011100000001011001: color_data = 8'b11111111;
		20'b00011100000001011010: color_data = 8'b11111111;
		20'b00011100000001011011: color_data = 8'b11111111;
		20'b00011100000001011100: color_data = 8'b11111111;
		20'b00011100000001011101: color_data = 8'b11111111;
		20'b00011100000001011110: color_data = 8'b11111111;
		20'b00011100000001011111: color_data = 8'b10010010;
		20'b00011100000001101000: color_data = 8'b10010010;
		20'b00011100000001101001: color_data = 8'b11111111;
		20'b00011100000001101010: color_data = 8'b11111111;
		20'b00011100000001101011: color_data = 8'b11111111;
		20'b00011100000001101100: color_data = 8'b11111111;
		20'b00011100000001101101: color_data = 8'b11111111;
		20'b00011100000001101110: color_data = 8'b11111111;
		20'b00011100000001101111: color_data = 8'b11111111;
		20'b00011100000001110000: color_data = 8'b11111111;
		20'b00011100000001110001: color_data = 8'b11111111;
		20'b00011100000001110010: color_data = 8'b10010010;
		20'b00011100000010000101: color_data = 8'b11011011;
		20'b00011100000010000110: color_data = 8'b11111111;
		20'b00011100000010000111: color_data = 8'b11111111;
		20'b00011100000010001000: color_data = 8'b11111111;
		20'b00011100000010001001: color_data = 8'b11111111;
		20'b00011100000010001010: color_data = 8'b11111111;
		20'b00011100000010001011: color_data = 8'b11111111;
		20'b00011100000010001100: color_data = 8'b11111111;
		20'b00011100000010001101: color_data = 8'b11111111;
		20'b00011100000010001110: color_data = 8'b11111111;
		20'b00011100000010011000: color_data = 8'b11011011;
		20'b00011100000010011001: color_data = 8'b11111111;
		20'b00011100000010011010: color_data = 8'b11111111;
		20'b00011100000010011011: color_data = 8'b11111111;
		20'b00011100000010011100: color_data = 8'b11111111;
		20'b00011100000010011101: color_data = 8'b11111111;
		20'b00011100000010011110: color_data = 8'b11111111;
		20'b00011100000010011111: color_data = 8'b11111111;
		20'b00011100000010100000: color_data = 8'b11111111;
		20'b00011100000010100001: color_data = 8'b11011011;
		20'b00011100000010110100: color_data = 8'b10010010;
		20'b00011100000010110101: color_data = 8'b11111111;
		20'b00011100000010110110: color_data = 8'b11111111;
		20'b00011100000010110111: color_data = 8'b11111111;
		20'b00011100000010111000: color_data = 8'b11111111;
		20'b00011100000010111001: color_data = 8'b11111111;
		20'b00011100000010111010: color_data = 8'b11111111;
		20'b00011100000010111011: color_data = 8'b11111111;
		20'b00011100000010111100: color_data = 8'b11111111;
		20'b00011100000010111101: color_data = 8'b11111111;
		20'b00011100000010111110: color_data = 8'b11011011;

		20'b00011100010000001001: color_data = 8'b11011011;
		20'b00011100010000001010: color_data = 8'b11111111;
		20'b00011100010000001011: color_data = 8'b11111111;
		20'b00011100010000001100: color_data = 8'b11111111;
		20'b00011100010000001101: color_data = 8'b11111111;
		20'b00011100010000001110: color_data = 8'b11111111;
		20'b00011100010000001111: color_data = 8'b11111111;
		20'b00011100010000010000: color_data = 8'b11111111;
		20'b00011100010000010001: color_data = 8'b11111111;
		20'b00011100010000010010: color_data = 8'b11111111;
		20'b00011100010000010011: color_data = 8'b10010010;
		20'b00011100010000111001: color_data = 8'b11111111;
		20'b00011100010000111010: color_data = 8'b11111111;
		20'b00011100010000111011: color_data = 8'b11111111;
		20'b00011100010000111100: color_data = 8'b11111111;
		20'b00011100010000111101: color_data = 8'b11111111;
		20'b00011100010000111110: color_data = 8'b11111111;
		20'b00011100010000111111: color_data = 8'b11111111;
		20'b00011100010001000000: color_data = 8'b11111111;
		20'b00011100010001000001: color_data = 8'b11111111;
		20'b00011100010001000010: color_data = 8'b11011011;
		20'b00011100010001010101: color_data = 8'b10010010;
		20'b00011100010001010110: color_data = 8'b11111111;
		20'b00011100010001010111: color_data = 8'b11111111;
		20'b00011100010001011000: color_data = 8'b11111111;
		20'b00011100010001011001: color_data = 8'b11111111;
		20'b00011100010001011010: color_data = 8'b11111111;
		20'b00011100010001011011: color_data = 8'b11111111;
		20'b00011100010001011100: color_data = 8'b11111111;
		20'b00011100010001011101: color_data = 8'b11111111;
		20'b00011100010001011110: color_data = 8'b11111111;
		20'b00011100010001011111: color_data = 8'b10010010;
		20'b00011100010001101000: color_data = 8'b10010010;
		20'b00011100010001101001: color_data = 8'b11111111;
		20'b00011100010001101010: color_data = 8'b11111111;
		20'b00011100010001101011: color_data = 8'b11111111;
		20'b00011100010001101100: color_data = 8'b11111111;
		20'b00011100010001101101: color_data = 8'b11111111;
		20'b00011100010001101110: color_data = 8'b11111111;
		20'b00011100010001101111: color_data = 8'b11111111;
		20'b00011100010001110000: color_data = 8'b11111111;
		20'b00011100010001110001: color_data = 8'b11111111;
		20'b00011100010001110010: color_data = 8'b10010010;
		20'b00011100010010000101: color_data = 8'b11011011;
		20'b00011100010010000110: color_data = 8'b11111111;
		20'b00011100010010000111: color_data = 8'b11111111;
		20'b00011100010010001000: color_data = 8'b11111111;
		20'b00011100010010001001: color_data = 8'b11111111;
		20'b00011100010010001010: color_data = 8'b11111111;
		20'b00011100010010001011: color_data = 8'b11111111;
		20'b00011100010010001100: color_data = 8'b11111111;
		20'b00011100010010001101: color_data = 8'b11111111;
		20'b00011100010010001110: color_data = 8'b11111111;
		20'b00011100010010011000: color_data = 8'b11011011;
		20'b00011100010010011001: color_data = 8'b11111111;
		20'b00011100010010011010: color_data = 8'b11111111;
		20'b00011100010010011011: color_data = 8'b11111111;
		20'b00011100010010011100: color_data = 8'b11111111;
		20'b00011100010010011101: color_data = 8'b11111111;
		20'b00011100010010011110: color_data = 8'b11111111;
		20'b00011100010010011111: color_data = 8'b11111111;
		20'b00011100010010100000: color_data = 8'b11111111;
		20'b00011100010010100001: color_data = 8'b11011011;
		20'b00011100010010110100: color_data = 8'b10010010;
		20'b00011100010010110101: color_data = 8'b11111111;
		20'b00011100010010110110: color_data = 8'b11111111;
		20'b00011100010010110111: color_data = 8'b11111111;
		20'b00011100010010111000: color_data = 8'b11111111;
		20'b00011100010010111001: color_data = 8'b11111111;
		20'b00011100010010111010: color_data = 8'b11111111;
		20'b00011100010010111011: color_data = 8'b11111111;
		20'b00011100010010111100: color_data = 8'b11111111;
		20'b00011100010010111101: color_data = 8'b11111111;
		20'b00011100010010111110: color_data = 8'b11011011;

		20'b00011100100000001001: color_data = 8'b11011011;
		20'b00011100100000001010: color_data = 8'b11111111;
		20'b00011100100000001011: color_data = 8'b11111111;
		20'b00011100100000001100: color_data = 8'b11111111;
		20'b00011100100000001101: color_data = 8'b11111111;
		20'b00011100100000001110: color_data = 8'b11111111;
		20'b00011100100000001111: color_data = 8'b11111111;
		20'b00011100100000010000: color_data = 8'b11111111;
		20'b00011100100000010001: color_data = 8'b11111111;
		20'b00011100100000010010: color_data = 8'b11111111;
		20'b00011100100000010011: color_data = 8'b10010010;
		20'b00011100100000111001: color_data = 8'b11111111;
		20'b00011100100000111010: color_data = 8'b11111111;
		20'b00011100100000111011: color_data = 8'b11111111;
		20'b00011100100000111100: color_data = 8'b11111111;
		20'b00011100100000111101: color_data = 8'b11111111;
		20'b00011100100000111110: color_data = 8'b11111111;
		20'b00011100100000111111: color_data = 8'b11111111;
		20'b00011100100001000000: color_data = 8'b11111111;
		20'b00011100100001000001: color_data = 8'b11111111;
		20'b00011100100001000010: color_data = 8'b11111111;
		20'b00011100100001000011: color_data = 8'b11011011;
		20'b00011100100001000100: color_data = 8'b11011011;
		20'b00011100100001000101: color_data = 8'b11011011;
		20'b00011100100001000110: color_data = 8'b11011011;
		20'b00011100100001000111: color_data = 8'b11011011;
		20'b00011100100001001000: color_data = 8'b11011011;
		20'b00011100100001001001: color_data = 8'b11011011;
		20'b00011100100001001010: color_data = 8'b11011011;
		20'b00011100100001001011: color_data = 8'b11011011;
		20'b00011100100001001100: color_data = 8'b11011011;
		20'b00011100100001001101: color_data = 8'b11011011;
		20'b00011100100001001110: color_data = 8'b11011011;
		20'b00011100100001001111: color_data = 8'b11011011;
		20'b00011100100001010000: color_data = 8'b11011011;
		20'b00011100100001010001: color_data = 8'b11011011;
		20'b00011100100001010010: color_data = 8'b11011011;
		20'b00011100100001010011: color_data = 8'b11011011;
		20'b00011100100001010100: color_data = 8'b11011011;
		20'b00011100100001010101: color_data = 8'b11011011;
		20'b00011100100001010110: color_data = 8'b11111111;
		20'b00011100100001010111: color_data = 8'b11111111;
		20'b00011100100001011000: color_data = 8'b11111111;
		20'b00011100100001011001: color_data = 8'b11111111;
		20'b00011100100001011010: color_data = 8'b11111111;
		20'b00011100100001011011: color_data = 8'b11111111;
		20'b00011100100001011100: color_data = 8'b11111111;
		20'b00011100100001011101: color_data = 8'b11111111;
		20'b00011100100001011110: color_data = 8'b11111111;
		20'b00011100100001011111: color_data = 8'b10010010;
		20'b00011100100001101000: color_data = 8'b10010010;
		20'b00011100100001101001: color_data = 8'b11111111;
		20'b00011100100001101010: color_data = 8'b11111111;
		20'b00011100100001101011: color_data = 8'b11111111;
		20'b00011100100001101100: color_data = 8'b11111111;
		20'b00011100100001101101: color_data = 8'b11111111;
		20'b00011100100001101110: color_data = 8'b11111111;
		20'b00011100100001101111: color_data = 8'b11111111;
		20'b00011100100001110000: color_data = 8'b11111111;
		20'b00011100100001110001: color_data = 8'b11111111;
		20'b00011100100001110010: color_data = 8'b10010010;
		20'b00011100100010000101: color_data = 8'b11011011;
		20'b00011100100010000110: color_data = 8'b11111111;
		20'b00011100100010000111: color_data = 8'b11111111;
		20'b00011100100010001000: color_data = 8'b11111111;
		20'b00011100100010001001: color_data = 8'b11111111;
		20'b00011100100010001010: color_data = 8'b11111111;
		20'b00011100100010001011: color_data = 8'b11111111;
		20'b00011100100010001100: color_data = 8'b11111111;
		20'b00011100100010001101: color_data = 8'b11111111;
		20'b00011100100010001110: color_data = 8'b11111111;
		20'b00011100100010011000: color_data = 8'b11011011;
		20'b00011100100010011001: color_data = 8'b11111111;
		20'b00011100100010011010: color_data = 8'b11111111;
		20'b00011100100010011011: color_data = 8'b11111111;
		20'b00011100100010011100: color_data = 8'b11111111;
		20'b00011100100010011101: color_data = 8'b11111111;
		20'b00011100100010011110: color_data = 8'b11111111;
		20'b00011100100010011111: color_data = 8'b11111111;
		20'b00011100100010100000: color_data = 8'b11111111;
		20'b00011100100010100001: color_data = 8'b11111111;
		20'b00011100100010100010: color_data = 8'b10010010;
		20'b00011100100010100011: color_data = 8'b11011011;
		20'b00011100100010100100: color_data = 8'b11011011;
		20'b00011100100010100101: color_data = 8'b11011011;
		20'b00011100100010100110: color_data = 8'b11011011;
		20'b00011100100010100111: color_data = 8'b11011011;
		20'b00011100100010101000: color_data = 8'b11011011;
		20'b00011100100010101001: color_data = 8'b11011011;
		20'b00011100100010101010: color_data = 8'b11011011;
		20'b00011100100010101011: color_data = 8'b11011011;
		20'b00011100100010101100: color_data = 8'b11011011;
		20'b00011100100010101101: color_data = 8'b11011011;
		20'b00011100100010101110: color_data = 8'b11011011;
		20'b00011100100010101111: color_data = 8'b11011011;
		20'b00011100100010110000: color_data = 8'b11011011;
		20'b00011100100010110001: color_data = 8'b11011011;
		20'b00011100100010110010: color_data = 8'b11011011;
		20'b00011100100010110011: color_data = 8'b11011011;
		20'b00011100100010110100: color_data = 8'b11011011;
		20'b00011100100010110101: color_data = 8'b11111111;
		20'b00011100100010110110: color_data = 8'b11111111;
		20'b00011100100010110111: color_data = 8'b11111111;
		20'b00011100100010111000: color_data = 8'b11111111;
		20'b00011100100010111001: color_data = 8'b11111111;
		20'b00011100100010111010: color_data = 8'b11111111;
		20'b00011100100010111011: color_data = 8'b11111111;
		20'b00011100100010111100: color_data = 8'b11111111;
		20'b00011100100010111101: color_data = 8'b11111111;
		20'b00011100100010111110: color_data = 8'b11011011;

		20'b00011100110000001001: color_data = 8'b11011011;
		20'b00011100110000001010: color_data = 8'b11111111;
		20'b00011100110000001011: color_data = 8'b11111111;
		20'b00011100110000001100: color_data = 8'b11111111;
		20'b00011100110000001101: color_data = 8'b11111111;
		20'b00011100110000001110: color_data = 8'b11111111;
		20'b00011100110000001111: color_data = 8'b11111111;
		20'b00011100110000010000: color_data = 8'b11111111;
		20'b00011100110000010001: color_data = 8'b11111111;
		20'b00011100110000010010: color_data = 8'b11111111;
		20'b00011100110000010011: color_data = 8'b10010010;
		20'b00011100110000111001: color_data = 8'b11111111;
		20'b00011100110000111010: color_data = 8'b11111111;
		20'b00011100110000111011: color_data = 8'b11111111;
		20'b00011100110000111100: color_data = 8'b11111111;
		20'b00011100110000111101: color_data = 8'b11111111;
		20'b00011100110000111110: color_data = 8'b11111111;
		20'b00011100110000111111: color_data = 8'b11111111;
		20'b00011100110001000000: color_data = 8'b11111111;
		20'b00011100110001000001: color_data = 8'b11111111;
		20'b00011100110001000010: color_data = 8'b11111111;
		20'b00011100110001000011: color_data = 8'b11111111;
		20'b00011100110001000100: color_data = 8'b11111111;
		20'b00011100110001000101: color_data = 8'b11111111;
		20'b00011100110001000110: color_data = 8'b11111111;
		20'b00011100110001000111: color_data = 8'b11111111;
		20'b00011100110001001000: color_data = 8'b11111111;
		20'b00011100110001001001: color_data = 8'b11111111;
		20'b00011100110001001010: color_data = 8'b11111111;
		20'b00011100110001001011: color_data = 8'b11111111;
		20'b00011100110001001100: color_data = 8'b11111111;
		20'b00011100110001001101: color_data = 8'b11111111;
		20'b00011100110001001110: color_data = 8'b11111111;
		20'b00011100110001001111: color_data = 8'b11111111;
		20'b00011100110001010000: color_data = 8'b11111111;
		20'b00011100110001010001: color_data = 8'b11111111;
		20'b00011100110001010010: color_data = 8'b11111111;
		20'b00011100110001010011: color_data = 8'b11111111;
		20'b00011100110001010100: color_data = 8'b11111111;
		20'b00011100110001010101: color_data = 8'b11111111;
		20'b00011100110001010110: color_data = 8'b11111111;
		20'b00011100110001010111: color_data = 8'b11111111;
		20'b00011100110001011000: color_data = 8'b11111111;
		20'b00011100110001011001: color_data = 8'b11111111;
		20'b00011100110001011010: color_data = 8'b11111111;
		20'b00011100110001011011: color_data = 8'b11111111;
		20'b00011100110001011100: color_data = 8'b11111111;
		20'b00011100110001011101: color_data = 8'b11111111;
		20'b00011100110001011110: color_data = 8'b11111111;
		20'b00011100110001011111: color_data = 8'b10010010;
		20'b00011100110001101000: color_data = 8'b10010010;
		20'b00011100110001101001: color_data = 8'b11111111;
		20'b00011100110001101010: color_data = 8'b11111111;
		20'b00011100110001101011: color_data = 8'b11111111;
		20'b00011100110001101100: color_data = 8'b11111111;
		20'b00011100110001101101: color_data = 8'b11111111;
		20'b00011100110001101110: color_data = 8'b11111111;
		20'b00011100110001101111: color_data = 8'b11111111;
		20'b00011100110001110000: color_data = 8'b11111111;
		20'b00011100110001110001: color_data = 8'b11111111;
		20'b00011100110001110010: color_data = 8'b10010010;
		20'b00011100110010000101: color_data = 8'b11011011;
		20'b00011100110010000110: color_data = 8'b11111111;
		20'b00011100110010000111: color_data = 8'b11111111;
		20'b00011100110010001000: color_data = 8'b11111111;
		20'b00011100110010001001: color_data = 8'b11111111;
		20'b00011100110010001010: color_data = 8'b11111111;
		20'b00011100110010001011: color_data = 8'b11111111;
		20'b00011100110010001100: color_data = 8'b11111111;
		20'b00011100110010001101: color_data = 8'b11111111;
		20'b00011100110010001110: color_data = 8'b11111111;
		20'b00011100110010011000: color_data = 8'b11011011;
		20'b00011100110010011001: color_data = 8'b11111111;
		20'b00011100110010011010: color_data = 8'b11111111;
		20'b00011100110010011011: color_data = 8'b11111111;
		20'b00011100110010011100: color_data = 8'b11111111;
		20'b00011100110010011101: color_data = 8'b11111111;
		20'b00011100110010011110: color_data = 8'b11111111;
		20'b00011100110010011111: color_data = 8'b11111111;
		20'b00011100110010100000: color_data = 8'b11111111;
		20'b00011100110010100001: color_data = 8'b11111111;
		20'b00011100110010100010: color_data = 8'b11111111;
		20'b00011100110010100011: color_data = 8'b11111111;
		20'b00011100110010100100: color_data = 8'b11111111;
		20'b00011100110010100101: color_data = 8'b11111111;
		20'b00011100110010100110: color_data = 8'b11111111;
		20'b00011100110010100111: color_data = 8'b11111111;
		20'b00011100110010101000: color_data = 8'b11111111;
		20'b00011100110010101001: color_data = 8'b11111111;
		20'b00011100110010101010: color_data = 8'b11111111;
		20'b00011100110010101011: color_data = 8'b11111111;
		20'b00011100110010101100: color_data = 8'b11111111;
		20'b00011100110010101101: color_data = 8'b11111111;
		20'b00011100110010101110: color_data = 8'b11111111;
		20'b00011100110010101111: color_data = 8'b11111111;
		20'b00011100110010110000: color_data = 8'b11111111;
		20'b00011100110010110001: color_data = 8'b11111111;
		20'b00011100110010110010: color_data = 8'b11111111;
		20'b00011100110010110011: color_data = 8'b11111111;
		20'b00011100110010110100: color_data = 8'b11111111;
		20'b00011100110010110101: color_data = 8'b11111111;
		20'b00011100110010110110: color_data = 8'b11111111;
		20'b00011100110010110111: color_data = 8'b11111111;
		20'b00011100110010111000: color_data = 8'b11111111;
		20'b00011100110010111001: color_data = 8'b11111111;
		20'b00011100110010111010: color_data = 8'b11111111;
		20'b00011100110010111011: color_data = 8'b11111111;
		20'b00011100110010111100: color_data = 8'b11111111;
		20'b00011100110010111101: color_data = 8'b11111111;
		20'b00011100110010111110: color_data = 8'b11011011;

		20'b00011101000000001001: color_data = 8'b11011011;
		20'b00011101000000001010: color_data = 8'b11111111;
		20'b00011101000000001011: color_data = 8'b11111111;
		20'b00011101000000001100: color_data = 8'b11111111;
		20'b00011101000000001101: color_data = 8'b11111111;
		20'b00011101000000001110: color_data = 8'b11111111;
		20'b00011101000000001111: color_data = 8'b11111111;
		20'b00011101000000010000: color_data = 8'b11111111;
		20'b00011101000000010001: color_data = 8'b11111111;
		20'b00011101000000010010: color_data = 8'b11111111;
		20'b00011101000000010011: color_data = 8'b10010010;
		20'b00011101000000111001: color_data = 8'b11111111;
		20'b00011101000000111010: color_data = 8'b11111111;
		20'b00011101000000111011: color_data = 8'b11111111;
		20'b00011101000000111100: color_data = 8'b11111111;
		20'b00011101000000111101: color_data = 8'b11111111;
		20'b00011101000000111110: color_data = 8'b11111111;
		20'b00011101000000111111: color_data = 8'b11111111;
		20'b00011101000001000000: color_data = 8'b11111111;
		20'b00011101000001000001: color_data = 8'b11111111;
		20'b00011101000001000010: color_data = 8'b11111111;
		20'b00011101000001000011: color_data = 8'b11111111;
		20'b00011101000001000100: color_data = 8'b11111111;
		20'b00011101000001000101: color_data = 8'b11111111;
		20'b00011101000001000110: color_data = 8'b11111111;
		20'b00011101000001000111: color_data = 8'b11111111;
		20'b00011101000001001000: color_data = 8'b11111111;
		20'b00011101000001001001: color_data = 8'b11111111;
		20'b00011101000001001010: color_data = 8'b11111111;
		20'b00011101000001001011: color_data = 8'b11111111;
		20'b00011101000001001100: color_data = 8'b11111111;
		20'b00011101000001001101: color_data = 8'b11111111;
		20'b00011101000001001110: color_data = 8'b11111111;
		20'b00011101000001001111: color_data = 8'b11111111;
		20'b00011101000001010000: color_data = 8'b11111111;
		20'b00011101000001010001: color_data = 8'b11111111;
		20'b00011101000001010010: color_data = 8'b11111111;
		20'b00011101000001010011: color_data = 8'b11111111;
		20'b00011101000001010100: color_data = 8'b11111111;
		20'b00011101000001010101: color_data = 8'b11111111;
		20'b00011101000001010110: color_data = 8'b11111111;
		20'b00011101000001010111: color_data = 8'b11111111;
		20'b00011101000001011000: color_data = 8'b11111111;
		20'b00011101000001011001: color_data = 8'b11111111;
		20'b00011101000001011010: color_data = 8'b11111111;
		20'b00011101000001011011: color_data = 8'b11111111;
		20'b00011101000001011100: color_data = 8'b11111111;
		20'b00011101000001011101: color_data = 8'b11111111;
		20'b00011101000001011110: color_data = 8'b11111111;
		20'b00011101000001011111: color_data = 8'b10010010;
		20'b00011101000001101000: color_data = 8'b10010010;
		20'b00011101000001101001: color_data = 8'b11111111;
		20'b00011101000001101010: color_data = 8'b11111111;
		20'b00011101000001101011: color_data = 8'b11111111;
		20'b00011101000001101100: color_data = 8'b11111111;
		20'b00011101000001101101: color_data = 8'b11111111;
		20'b00011101000001101110: color_data = 8'b11111111;
		20'b00011101000001101111: color_data = 8'b11111111;
		20'b00011101000001110000: color_data = 8'b11111111;
		20'b00011101000001110001: color_data = 8'b11111111;
		20'b00011101000001110010: color_data = 8'b10010010;
		20'b00011101000010000101: color_data = 8'b11011011;
		20'b00011101000010000110: color_data = 8'b11111111;
		20'b00011101000010000111: color_data = 8'b11111111;
		20'b00011101000010001000: color_data = 8'b11111111;
		20'b00011101000010001001: color_data = 8'b11111111;
		20'b00011101000010001010: color_data = 8'b11111111;
		20'b00011101000010001011: color_data = 8'b11111111;
		20'b00011101000010001100: color_data = 8'b11111111;
		20'b00011101000010001101: color_data = 8'b11111111;
		20'b00011101000010001110: color_data = 8'b11111111;
		20'b00011101000010011000: color_data = 8'b11011011;
		20'b00011101000010011001: color_data = 8'b11111111;
		20'b00011101000010011010: color_data = 8'b11111111;
		20'b00011101000010011011: color_data = 8'b11111111;
		20'b00011101000010011100: color_data = 8'b11111111;
		20'b00011101000010011101: color_data = 8'b11111111;
		20'b00011101000010011110: color_data = 8'b11111111;
		20'b00011101000010011111: color_data = 8'b11111111;
		20'b00011101000010100000: color_data = 8'b11111111;
		20'b00011101000010100001: color_data = 8'b11111111;
		20'b00011101000010100010: color_data = 8'b11111111;
		20'b00011101000010100011: color_data = 8'b11111111;
		20'b00011101000010100100: color_data = 8'b11111111;
		20'b00011101000010100101: color_data = 8'b11111111;
		20'b00011101000010100110: color_data = 8'b11111111;
		20'b00011101000010100111: color_data = 8'b11111111;
		20'b00011101000010101000: color_data = 8'b11111111;
		20'b00011101000010101001: color_data = 8'b11111111;
		20'b00011101000010101010: color_data = 8'b11111111;
		20'b00011101000010101011: color_data = 8'b11111111;
		20'b00011101000010101100: color_data = 8'b11111111;
		20'b00011101000010101101: color_data = 8'b11111111;
		20'b00011101000010101110: color_data = 8'b11111111;
		20'b00011101000010101111: color_data = 8'b11111111;
		20'b00011101000010110000: color_data = 8'b11111111;
		20'b00011101000010110001: color_data = 8'b11111111;
		20'b00011101000010110010: color_data = 8'b11111111;
		20'b00011101000010110011: color_data = 8'b11111111;
		20'b00011101000010110100: color_data = 8'b11111111;
		20'b00011101000010110101: color_data = 8'b11111111;
		20'b00011101000010110110: color_data = 8'b11111111;
		20'b00011101000010110111: color_data = 8'b11111111;
		20'b00011101000010111000: color_data = 8'b11111111;
		20'b00011101000010111001: color_data = 8'b11111111;
		20'b00011101000010111010: color_data = 8'b11111111;
		20'b00011101000010111011: color_data = 8'b11111111;
		20'b00011101000010111100: color_data = 8'b11111111;
		20'b00011101000010111101: color_data = 8'b11111111;
		20'b00011101000010111110: color_data = 8'b11011011;

		20'b00011101010000001001: color_data = 8'b11011011;
		20'b00011101010000001010: color_data = 8'b11111111;
		20'b00011101010000001011: color_data = 8'b11111111;
		20'b00011101010000001100: color_data = 8'b11111111;
		20'b00011101010000001101: color_data = 8'b11111111;
		20'b00011101010000001110: color_data = 8'b11111111;
		20'b00011101010000001111: color_data = 8'b11111111;
		20'b00011101010000010000: color_data = 8'b11111111;
		20'b00011101010000010001: color_data = 8'b11111111;
		20'b00011101010000010010: color_data = 8'b11111111;
		20'b00011101010000010011: color_data = 8'b10010010;
		20'b00011101010000111001: color_data = 8'b11111111;
		20'b00011101010000111010: color_data = 8'b11111111;
		20'b00011101010000111011: color_data = 8'b11111111;
		20'b00011101010000111100: color_data = 8'b11111111;
		20'b00011101010000111101: color_data = 8'b11111111;
		20'b00011101010000111110: color_data = 8'b11111111;
		20'b00011101010000111111: color_data = 8'b11111111;
		20'b00011101010001000000: color_data = 8'b11111111;
		20'b00011101010001000001: color_data = 8'b11111111;
		20'b00011101010001000010: color_data = 8'b11111111;
		20'b00011101010001000011: color_data = 8'b11111111;
		20'b00011101010001000100: color_data = 8'b11111111;
		20'b00011101010001000101: color_data = 8'b11111111;
		20'b00011101010001000110: color_data = 8'b11111111;
		20'b00011101010001000111: color_data = 8'b11111111;
		20'b00011101010001001000: color_data = 8'b11111111;
		20'b00011101010001001001: color_data = 8'b11111111;
		20'b00011101010001001010: color_data = 8'b11111111;
		20'b00011101010001001011: color_data = 8'b11111111;
		20'b00011101010001001100: color_data = 8'b11111111;
		20'b00011101010001001101: color_data = 8'b11111111;
		20'b00011101010001001110: color_data = 8'b11111111;
		20'b00011101010001001111: color_data = 8'b11111111;
		20'b00011101010001010000: color_data = 8'b11111111;
		20'b00011101010001010001: color_data = 8'b11111111;
		20'b00011101010001010010: color_data = 8'b11111111;
		20'b00011101010001010011: color_data = 8'b11111111;
		20'b00011101010001010100: color_data = 8'b11111111;
		20'b00011101010001010101: color_data = 8'b11111111;
		20'b00011101010001010110: color_data = 8'b11111111;
		20'b00011101010001010111: color_data = 8'b11111111;
		20'b00011101010001011000: color_data = 8'b11111111;
		20'b00011101010001011001: color_data = 8'b11111111;
		20'b00011101010001011010: color_data = 8'b11111111;
		20'b00011101010001011011: color_data = 8'b11111111;
		20'b00011101010001011100: color_data = 8'b11111111;
		20'b00011101010001011101: color_data = 8'b11111111;
		20'b00011101010001011110: color_data = 8'b11111111;
		20'b00011101010001011111: color_data = 8'b10010010;
		20'b00011101010001101000: color_data = 8'b10010010;
		20'b00011101010001101001: color_data = 8'b11111111;
		20'b00011101010001101010: color_data = 8'b11111111;
		20'b00011101010001101011: color_data = 8'b11111111;
		20'b00011101010001101100: color_data = 8'b11111111;
		20'b00011101010001101101: color_data = 8'b11111111;
		20'b00011101010001101110: color_data = 8'b11111111;
		20'b00011101010001101111: color_data = 8'b11111111;
		20'b00011101010001110000: color_data = 8'b11111111;
		20'b00011101010001110001: color_data = 8'b11111111;
		20'b00011101010001110010: color_data = 8'b10010010;
		20'b00011101010010000101: color_data = 8'b11011011;
		20'b00011101010010000110: color_data = 8'b11111111;
		20'b00011101010010000111: color_data = 8'b11111111;
		20'b00011101010010001000: color_data = 8'b11111111;
		20'b00011101010010001001: color_data = 8'b11111111;
		20'b00011101010010001010: color_data = 8'b11111111;
		20'b00011101010010001011: color_data = 8'b11111111;
		20'b00011101010010001100: color_data = 8'b11111111;
		20'b00011101010010001101: color_data = 8'b11111111;
		20'b00011101010010001110: color_data = 8'b11111111;
		20'b00011101010010011000: color_data = 8'b11011011;
		20'b00011101010010011001: color_data = 8'b11111111;
		20'b00011101010010011010: color_data = 8'b11111111;
		20'b00011101010010011011: color_data = 8'b11111111;
		20'b00011101010010011100: color_data = 8'b11111111;
		20'b00011101010010011101: color_data = 8'b11111111;
		20'b00011101010010011110: color_data = 8'b11111111;
		20'b00011101010010011111: color_data = 8'b11111111;
		20'b00011101010010100000: color_data = 8'b11111111;
		20'b00011101010010100001: color_data = 8'b11111111;
		20'b00011101010010100010: color_data = 8'b11111111;
		20'b00011101010010100011: color_data = 8'b11111111;
		20'b00011101010010100100: color_data = 8'b11111111;
		20'b00011101010010100101: color_data = 8'b11111111;
		20'b00011101010010100110: color_data = 8'b11111111;
		20'b00011101010010100111: color_data = 8'b11111111;
		20'b00011101010010101000: color_data = 8'b11111111;
		20'b00011101010010101001: color_data = 8'b11111111;
		20'b00011101010010101010: color_data = 8'b11111111;
		20'b00011101010010101011: color_data = 8'b11111111;
		20'b00011101010010101100: color_data = 8'b11111111;
		20'b00011101010010101101: color_data = 8'b11111111;
		20'b00011101010010101110: color_data = 8'b11111111;
		20'b00011101010010101111: color_data = 8'b11111111;
		20'b00011101010010110000: color_data = 8'b11111111;
		20'b00011101010010110001: color_data = 8'b11111111;
		20'b00011101010010110010: color_data = 8'b11111111;
		20'b00011101010010110011: color_data = 8'b11111111;
		20'b00011101010010110100: color_data = 8'b11111111;
		20'b00011101010010110101: color_data = 8'b11111111;
		20'b00011101010010110110: color_data = 8'b11111111;
		20'b00011101010010110111: color_data = 8'b11111111;
		20'b00011101010010111000: color_data = 8'b11111111;
		20'b00011101010010111001: color_data = 8'b11111111;
		20'b00011101010010111010: color_data = 8'b11111111;
		20'b00011101010010111011: color_data = 8'b11111111;
		20'b00011101010010111100: color_data = 8'b11111111;
		20'b00011101010010111101: color_data = 8'b11111111;
		20'b00011101010010111110: color_data = 8'b11011011;

		20'b00011101100000001001: color_data = 8'b11011011;
		20'b00011101100000001010: color_data = 8'b11111111;
		20'b00011101100000001011: color_data = 8'b11111111;
		20'b00011101100000001100: color_data = 8'b11111111;
		20'b00011101100000001101: color_data = 8'b11111111;
		20'b00011101100000001110: color_data = 8'b11111111;
		20'b00011101100000001111: color_data = 8'b11111111;
		20'b00011101100000010000: color_data = 8'b11111111;
		20'b00011101100000010001: color_data = 8'b11111111;
		20'b00011101100000010010: color_data = 8'b11111111;
		20'b00011101100000010011: color_data = 8'b10010010;
		20'b00011101100000111001: color_data = 8'b11111111;
		20'b00011101100000111010: color_data = 8'b11111111;
		20'b00011101100000111011: color_data = 8'b11111111;
		20'b00011101100000111100: color_data = 8'b11111111;
		20'b00011101100000111101: color_data = 8'b11111111;
		20'b00011101100000111110: color_data = 8'b11111111;
		20'b00011101100000111111: color_data = 8'b11111111;
		20'b00011101100001000000: color_data = 8'b11111111;
		20'b00011101100001000001: color_data = 8'b11111111;
		20'b00011101100001000010: color_data = 8'b11111111;
		20'b00011101100001000011: color_data = 8'b11111111;
		20'b00011101100001000100: color_data = 8'b11111111;
		20'b00011101100001000101: color_data = 8'b11111111;
		20'b00011101100001000110: color_data = 8'b11111111;
		20'b00011101100001000111: color_data = 8'b11111111;
		20'b00011101100001001000: color_data = 8'b11111111;
		20'b00011101100001001001: color_data = 8'b11111111;
		20'b00011101100001001010: color_data = 8'b11111111;
		20'b00011101100001001011: color_data = 8'b11111111;
		20'b00011101100001001100: color_data = 8'b11111111;
		20'b00011101100001001101: color_data = 8'b11111111;
		20'b00011101100001001110: color_data = 8'b11111111;
		20'b00011101100001001111: color_data = 8'b11111111;
		20'b00011101100001010000: color_data = 8'b11111111;
		20'b00011101100001010001: color_data = 8'b11111111;
		20'b00011101100001010010: color_data = 8'b11111111;
		20'b00011101100001010011: color_data = 8'b11111111;
		20'b00011101100001010100: color_data = 8'b11111111;
		20'b00011101100001010101: color_data = 8'b11111111;
		20'b00011101100001010110: color_data = 8'b11111111;
		20'b00011101100001010111: color_data = 8'b11111111;
		20'b00011101100001011000: color_data = 8'b11111111;
		20'b00011101100001011001: color_data = 8'b11111111;
		20'b00011101100001011010: color_data = 8'b11111111;
		20'b00011101100001011011: color_data = 8'b11111111;
		20'b00011101100001011100: color_data = 8'b11111111;
		20'b00011101100001011101: color_data = 8'b11111111;
		20'b00011101100001011110: color_data = 8'b11111111;
		20'b00011101100001011111: color_data = 8'b10010010;
		20'b00011101100001101000: color_data = 8'b10010010;
		20'b00011101100001101001: color_data = 8'b11111111;
		20'b00011101100001101010: color_data = 8'b11111111;
		20'b00011101100001101011: color_data = 8'b11111111;
		20'b00011101100001101100: color_data = 8'b11111111;
		20'b00011101100001101101: color_data = 8'b11111111;
		20'b00011101100001101110: color_data = 8'b11111111;
		20'b00011101100001101111: color_data = 8'b11111111;
		20'b00011101100001110000: color_data = 8'b11111111;
		20'b00011101100001110001: color_data = 8'b11111111;
		20'b00011101100001110010: color_data = 8'b10010010;
		20'b00011101100010000101: color_data = 8'b11011011;
		20'b00011101100010000110: color_data = 8'b11111111;
		20'b00011101100010000111: color_data = 8'b11111111;
		20'b00011101100010001000: color_data = 8'b11111111;
		20'b00011101100010001001: color_data = 8'b11111111;
		20'b00011101100010001010: color_data = 8'b11111111;
		20'b00011101100010001011: color_data = 8'b11111111;
		20'b00011101100010001100: color_data = 8'b11111111;
		20'b00011101100010001101: color_data = 8'b11111111;
		20'b00011101100010001110: color_data = 8'b11111111;
		20'b00011101100010011000: color_data = 8'b11011011;
		20'b00011101100010011001: color_data = 8'b11111111;
		20'b00011101100010011010: color_data = 8'b11111111;
		20'b00011101100010011011: color_data = 8'b11111111;
		20'b00011101100010011100: color_data = 8'b11111111;
		20'b00011101100010011101: color_data = 8'b11111111;
		20'b00011101100010011110: color_data = 8'b11111111;
		20'b00011101100010011111: color_data = 8'b11111111;
		20'b00011101100010100000: color_data = 8'b11111111;
		20'b00011101100010100001: color_data = 8'b11111111;
		20'b00011101100010100010: color_data = 8'b11111111;
		20'b00011101100010100011: color_data = 8'b11111111;
		20'b00011101100010100100: color_data = 8'b11111111;
		20'b00011101100010100101: color_data = 8'b11111111;
		20'b00011101100010100110: color_data = 8'b11111111;
		20'b00011101100010100111: color_data = 8'b11111111;
		20'b00011101100010101000: color_data = 8'b11111111;
		20'b00011101100010101001: color_data = 8'b11111111;
		20'b00011101100010101010: color_data = 8'b11111111;
		20'b00011101100010101011: color_data = 8'b11111111;
		20'b00011101100010101100: color_data = 8'b11111111;
		20'b00011101100010101101: color_data = 8'b11111111;
		20'b00011101100010101110: color_data = 8'b11111111;
		20'b00011101100010101111: color_data = 8'b11111111;
		20'b00011101100010110000: color_data = 8'b11111111;
		20'b00011101100010110001: color_data = 8'b11111111;
		20'b00011101100010110010: color_data = 8'b11111111;
		20'b00011101100010110011: color_data = 8'b11111111;
		20'b00011101100010110100: color_data = 8'b11111111;
		20'b00011101100010110101: color_data = 8'b11111111;
		20'b00011101100010110110: color_data = 8'b11111111;
		20'b00011101100010110111: color_data = 8'b11111111;
		20'b00011101100010111000: color_data = 8'b11111111;
		20'b00011101100010111001: color_data = 8'b11111111;
		20'b00011101100010111010: color_data = 8'b11111111;
		20'b00011101100010111011: color_data = 8'b11111111;
		20'b00011101100010111100: color_data = 8'b11111111;
		20'b00011101100010111101: color_data = 8'b11111111;
		20'b00011101100010111110: color_data = 8'b11011011;

		20'b00011101110000001001: color_data = 8'b11011011;
		20'b00011101110000001010: color_data = 8'b11111111;
		20'b00011101110000001011: color_data = 8'b11111111;
		20'b00011101110000001100: color_data = 8'b11111111;
		20'b00011101110000001101: color_data = 8'b11111111;
		20'b00011101110000001110: color_data = 8'b11111111;
		20'b00011101110000001111: color_data = 8'b11111111;
		20'b00011101110000010000: color_data = 8'b11111111;
		20'b00011101110000010001: color_data = 8'b11111111;
		20'b00011101110000010010: color_data = 8'b11111111;
		20'b00011101110000010011: color_data = 8'b10010010;
		20'b00011101110000111001: color_data = 8'b11111111;
		20'b00011101110000111010: color_data = 8'b11111111;
		20'b00011101110000111011: color_data = 8'b11111111;
		20'b00011101110000111100: color_data = 8'b11111111;
		20'b00011101110000111101: color_data = 8'b11111111;
		20'b00011101110000111110: color_data = 8'b11111111;
		20'b00011101110000111111: color_data = 8'b11111111;
		20'b00011101110001000000: color_data = 8'b11111111;
		20'b00011101110001000001: color_data = 8'b11111111;
		20'b00011101110001000010: color_data = 8'b11111111;
		20'b00011101110001000011: color_data = 8'b11111111;
		20'b00011101110001000100: color_data = 8'b11111111;
		20'b00011101110001000101: color_data = 8'b11111111;
		20'b00011101110001000110: color_data = 8'b11111111;
		20'b00011101110001000111: color_data = 8'b11111111;
		20'b00011101110001001000: color_data = 8'b11111111;
		20'b00011101110001001001: color_data = 8'b11111111;
		20'b00011101110001001010: color_data = 8'b11111111;
		20'b00011101110001001011: color_data = 8'b11111111;
		20'b00011101110001001100: color_data = 8'b11111111;
		20'b00011101110001001101: color_data = 8'b11111111;
		20'b00011101110001001110: color_data = 8'b11111111;
		20'b00011101110001001111: color_data = 8'b11111111;
		20'b00011101110001010000: color_data = 8'b11111111;
		20'b00011101110001010001: color_data = 8'b11111111;
		20'b00011101110001010010: color_data = 8'b11111111;
		20'b00011101110001010011: color_data = 8'b11111111;
		20'b00011101110001010100: color_data = 8'b11111111;
		20'b00011101110001010101: color_data = 8'b11111111;
		20'b00011101110001010110: color_data = 8'b11111111;
		20'b00011101110001010111: color_data = 8'b11111111;
		20'b00011101110001011000: color_data = 8'b11111111;
		20'b00011101110001011001: color_data = 8'b11111111;
		20'b00011101110001011010: color_data = 8'b11111111;
		20'b00011101110001011011: color_data = 8'b11111111;
		20'b00011101110001011100: color_data = 8'b11111111;
		20'b00011101110001011101: color_data = 8'b11111111;
		20'b00011101110001011110: color_data = 8'b11111111;
		20'b00011101110001011111: color_data = 8'b10010010;
		20'b00011101110001101000: color_data = 8'b10010010;
		20'b00011101110001101001: color_data = 8'b11111111;
		20'b00011101110001101010: color_data = 8'b11111111;
		20'b00011101110001101011: color_data = 8'b11111111;
		20'b00011101110001101100: color_data = 8'b11111111;
		20'b00011101110001101101: color_data = 8'b11111111;
		20'b00011101110001101110: color_data = 8'b11111111;
		20'b00011101110001101111: color_data = 8'b11111111;
		20'b00011101110001110000: color_data = 8'b11111111;
		20'b00011101110001110001: color_data = 8'b11111111;
		20'b00011101110001110010: color_data = 8'b10010010;
		20'b00011101110010000101: color_data = 8'b11011011;
		20'b00011101110010000110: color_data = 8'b11111111;
		20'b00011101110010000111: color_data = 8'b11111111;
		20'b00011101110010001000: color_data = 8'b11111111;
		20'b00011101110010001001: color_data = 8'b11111111;
		20'b00011101110010001010: color_data = 8'b11111111;
		20'b00011101110010001011: color_data = 8'b11111111;
		20'b00011101110010001100: color_data = 8'b11111111;
		20'b00011101110010001101: color_data = 8'b11111111;
		20'b00011101110010001110: color_data = 8'b11111111;
		20'b00011101110010011000: color_data = 8'b11011011;
		20'b00011101110010011001: color_data = 8'b11111111;
		20'b00011101110010011010: color_data = 8'b11111111;
		20'b00011101110010011011: color_data = 8'b11111111;
		20'b00011101110010011100: color_data = 8'b11111111;
		20'b00011101110010011101: color_data = 8'b11111111;
		20'b00011101110010011110: color_data = 8'b11111111;
		20'b00011101110010011111: color_data = 8'b11111111;
		20'b00011101110010100000: color_data = 8'b11111111;
		20'b00011101110010100001: color_data = 8'b11111111;
		20'b00011101110010100010: color_data = 8'b11111111;
		20'b00011101110010100011: color_data = 8'b11111111;
		20'b00011101110010100100: color_data = 8'b11111111;
		20'b00011101110010100101: color_data = 8'b11111111;
		20'b00011101110010100110: color_data = 8'b11111111;
		20'b00011101110010100111: color_data = 8'b11111111;
		20'b00011101110010101000: color_data = 8'b11111111;
		20'b00011101110010101001: color_data = 8'b11111111;
		20'b00011101110010101010: color_data = 8'b11111111;
		20'b00011101110010101011: color_data = 8'b11111111;
		20'b00011101110010101100: color_data = 8'b11111111;
		20'b00011101110010101101: color_data = 8'b11111111;
		20'b00011101110010101110: color_data = 8'b11111111;
		20'b00011101110010101111: color_data = 8'b11111111;
		20'b00011101110010110000: color_data = 8'b11111111;
		20'b00011101110010110001: color_data = 8'b11111111;
		20'b00011101110010110010: color_data = 8'b11111111;
		20'b00011101110010110011: color_data = 8'b11111111;
		20'b00011101110010110100: color_data = 8'b11111111;
		20'b00011101110010110101: color_data = 8'b11111111;
		20'b00011101110010110110: color_data = 8'b11111111;
		20'b00011101110010110111: color_data = 8'b11111111;
		20'b00011101110010111000: color_data = 8'b11111111;
		20'b00011101110010111001: color_data = 8'b11111111;
		20'b00011101110010111010: color_data = 8'b11111111;
		20'b00011101110010111011: color_data = 8'b11111111;
		20'b00011101110010111100: color_data = 8'b11111111;
		20'b00011101110010111101: color_data = 8'b11111111;
		20'b00011101110010111110: color_data = 8'b11011011;

		20'b00011110000000001001: color_data = 8'b11011011;
		20'b00011110000000001010: color_data = 8'b11111111;
		20'b00011110000000001011: color_data = 8'b11111111;
		20'b00011110000000001100: color_data = 8'b11111111;
		20'b00011110000000001101: color_data = 8'b11111111;
		20'b00011110000000001110: color_data = 8'b11111111;
		20'b00011110000000001111: color_data = 8'b11111111;
		20'b00011110000000010000: color_data = 8'b11111111;
		20'b00011110000000010001: color_data = 8'b11111111;
		20'b00011110000000010010: color_data = 8'b11111111;
		20'b00011110000000010011: color_data = 8'b10010010;
		20'b00011110000000111001: color_data = 8'b11111111;
		20'b00011110000000111010: color_data = 8'b11111111;
		20'b00011110000000111011: color_data = 8'b11111111;
		20'b00011110000000111100: color_data = 8'b11111111;
		20'b00011110000000111101: color_data = 8'b11111111;
		20'b00011110000000111110: color_data = 8'b11111111;
		20'b00011110000000111111: color_data = 8'b11111111;
		20'b00011110000001000000: color_data = 8'b11111111;
		20'b00011110000001000001: color_data = 8'b11111111;
		20'b00011110000001000010: color_data = 8'b11111111;
		20'b00011110000001000011: color_data = 8'b11111111;
		20'b00011110000001000100: color_data = 8'b11111111;
		20'b00011110000001000101: color_data = 8'b11111111;
		20'b00011110000001000110: color_data = 8'b11111111;
		20'b00011110000001000111: color_data = 8'b11111111;
		20'b00011110000001001000: color_data = 8'b11111111;
		20'b00011110000001001001: color_data = 8'b11111111;
		20'b00011110000001001010: color_data = 8'b11111111;
		20'b00011110000001001011: color_data = 8'b11111111;
		20'b00011110000001001100: color_data = 8'b11111111;
		20'b00011110000001001101: color_data = 8'b11111111;
		20'b00011110000001001110: color_data = 8'b11111111;
		20'b00011110000001001111: color_data = 8'b11111111;
		20'b00011110000001010000: color_data = 8'b11111111;
		20'b00011110000001010001: color_data = 8'b11111111;
		20'b00011110000001010010: color_data = 8'b11111111;
		20'b00011110000001010011: color_data = 8'b11111111;
		20'b00011110000001010100: color_data = 8'b11111111;
		20'b00011110000001010101: color_data = 8'b11111111;
		20'b00011110000001010110: color_data = 8'b11111111;
		20'b00011110000001010111: color_data = 8'b11111111;
		20'b00011110000001011000: color_data = 8'b11111111;
		20'b00011110000001011001: color_data = 8'b11111111;
		20'b00011110000001011010: color_data = 8'b11111111;
		20'b00011110000001011011: color_data = 8'b11111111;
		20'b00011110000001011100: color_data = 8'b11111111;
		20'b00011110000001011101: color_data = 8'b11111111;
		20'b00011110000001011110: color_data = 8'b11111111;
		20'b00011110000001011111: color_data = 8'b10010010;
		20'b00011110000001101000: color_data = 8'b10010010;
		20'b00011110000001101001: color_data = 8'b11111111;
		20'b00011110000001101010: color_data = 8'b11111111;
		20'b00011110000001101011: color_data = 8'b11111111;
		20'b00011110000001101100: color_data = 8'b11111111;
		20'b00011110000001101101: color_data = 8'b11111111;
		20'b00011110000001101110: color_data = 8'b11111111;
		20'b00011110000001101111: color_data = 8'b11111111;
		20'b00011110000001110000: color_data = 8'b11111111;
		20'b00011110000001110001: color_data = 8'b11111111;
		20'b00011110000001110010: color_data = 8'b10010010;
		20'b00011110000010000101: color_data = 8'b11011011;
		20'b00011110000010000110: color_data = 8'b11111111;
		20'b00011110000010000111: color_data = 8'b11111111;
		20'b00011110000010001000: color_data = 8'b11111111;
		20'b00011110000010001001: color_data = 8'b11111111;
		20'b00011110000010001010: color_data = 8'b11111111;
		20'b00011110000010001011: color_data = 8'b11111111;
		20'b00011110000010001100: color_data = 8'b11111111;
		20'b00011110000010001101: color_data = 8'b11111111;
		20'b00011110000010001110: color_data = 8'b11111111;
		20'b00011110000010011000: color_data = 8'b11011011;
		20'b00011110000010011001: color_data = 8'b11111111;
		20'b00011110000010011010: color_data = 8'b11111111;
		20'b00011110000010011011: color_data = 8'b11111111;
		20'b00011110000010011100: color_data = 8'b11111111;
		20'b00011110000010011101: color_data = 8'b11111111;
		20'b00011110000010011110: color_data = 8'b11111111;
		20'b00011110000010011111: color_data = 8'b11111111;
		20'b00011110000010100000: color_data = 8'b11111111;
		20'b00011110000010100001: color_data = 8'b11111111;
		20'b00011110000010100010: color_data = 8'b11111111;
		20'b00011110000010100011: color_data = 8'b11111111;
		20'b00011110000010100100: color_data = 8'b11111111;
		20'b00011110000010100101: color_data = 8'b11111111;
		20'b00011110000010100110: color_data = 8'b11111111;
		20'b00011110000010100111: color_data = 8'b11111111;
		20'b00011110000010101000: color_data = 8'b11111111;
		20'b00011110000010101001: color_data = 8'b11111111;
		20'b00011110000010101010: color_data = 8'b11111111;
		20'b00011110000010101011: color_data = 8'b11111111;
		20'b00011110000010101100: color_data = 8'b11111111;
		20'b00011110000010101101: color_data = 8'b11111111;
		20'b00011110000010101110: color_data = 8'b11111111;
		20'b00011110000010101111: color_data = 8'b11111111;
		20'b00011110000010110000: color_data = 8'b11111111;
		20'b00011110000010110001: color_data = 8'b11111111;
		20'b00011110000010110010: color_data = 8'b11111111;
		20'b00011110000010110011: color_data = 8'b11111111;
		20'b00011110000010110100: color_data = 8'b11111111;
		20'b00011110000010110101: color_data = 8'b11111111;
		20'b00011110000010110110: color_data = 8'b11111111;
		20'b00011110000010110111: color_data = 8'b11111111;
		20'b00011110000010111000: color_data = 8'b11111111;
		20'b00011110000010111001: color_data = 8'b11111111;
		20'b00011110000010111010: color_data = 8'b11111111;
		20'b00011110000010111011: color_data = 8'b11111111;
		20'b00011110000010111100: color_data = 8'b11111111;
		20'b00011110000010111101: color_data = 8'b11111111;
		20'b00011110000010111110: color_data = 8'b11011011;

		20'b00011110010000001001: color_data = 8'b11011011;
		20'b00011110010000001010: color_data = 8'b11111111;
		20'b00011110010000001011: color_data = 8'b11111111;
		20'b00011110010000001100: color_data = 8'b11111111;
		20'b00011110010000001101: color_data = 8'b11111111;
		20'b00011110010000001110: color_data = 8'b11111111;
		20'b00011110010000001111: color_data = 8'b11111111;
		20'b00011110010000010000: color_data = 8'b11111111;
		20'b00011110010000010001: color_data = 8'b11111111;
		20'b00011110010000010010: color_data = 8'b11111111;
		20'b00011110010000010011: color_data = 8'b10010010;
		20'b00011110010000111001: color_data = 8'b11111111;
		20'b00011110010000111010: color_data = 8'b11111111;
		20'b00011110010000111011: color_data = 8'b11111111;
		20'b00011110010000111100: color_data = 8'b11111111;
		20'b00011110010000111101: color_data = 8'b11111111;
		20'b00011110010000111110: color_data = 8'b11111111;
		20'b00011110010000111111: color_data = 8'b11111111;
		20'b00011110010001000000: color_data = 8'b11111111;
		20'b00011110010001000001: color_data = 8'b11111111;
		20'b00011110010001000010: color_data = 8'b11111111;
		20'b00011110010001000011: color_data = 8'b11111111;
		20'b00011110010001000100: color_data = 8'b11111111;
		20'b00011110010001000101: color_data = 8'b11111111;
		20'b00011110010001000110: color_data = 8'b11111111;
		20'b00011110010001000111: color_data = 8'b11111111;
		20'b00011110010001001000: color_data = 8'b11111111;
		20'b00011110010001001001: color_data = 8'b11111111;
		20'b00011110010001001010: color_data = 8'b11111111;
		20'b00011110010001001011: color_data = 8'b11111111;
		20'b00011110010001001100: color_data = 8'b11111111;
		20'b00011110010001001101: color_data = 8'b11111111;
		20'b00011110010001001110: color_data = 8'b11111111;
		20'b00011110010001001111: color_data = 8'b11111111;
		20'b00011110010001010000: color_data = 8'b11111111;
		20'b00011110010001010001: color_data = 8'b11111111;
		20'b00011110010001010010: color_data = 8'b11111111;
		20'b00011110010001010011: color_data = 8'b11111111;
		20'b00011110010001010100: color_data = 8'b11111111;
		20'b00011110010001010101: color_data = 8'b11111111;
		20'b00011110010001010110: color_data = 8'b11111111;
		20'b00011110010001010111: color_data = 8'b11111111;
		20'b00011110010001011000: color_data = 8'b11111111;
		20'b00011110010001011001: color_data = 8'b11111111;
		20'b00011110010001011010: color_data = 8'b11111111;
		20'b00011110010001011011: color_data = 8'b11111111;
		20'b00011110010001011100: color_data = 8'b11111111;
		20'b00011110010001011101: color_data = 8'b11111111;
		20'b00011110010001011110: color_data = 8'b11111111;
		20'b00011110010001011111: color_data = 8'b10010010;
		20'b00011110010001101000: color_data = 8'b10010010;
		20'b00011110010001101001: color_data = 8'b11111111;
		20'b00011110010001101010: color_data = 8'b11111111;
		20'b00011110010001101011: color_data = 8'b11111111;
		20'b00011110010001101100: color_data = 8'b11111111;
		20'b00011110010001101101: color_data = 8'b11111111;
		20'b00011110010001101110: color_data = 8'b11111111;
		20'b00011110010001101111: color_data = 8'b11111111;
		20'b00011110010001110000: color_data = 8'b11111111;
		20'b00011110010001110001: color_data = 8'b11111111;
		20'b00011110010001110010: color_data = 8'b10010010;
		20'b00011110010010000101: color_data = 8'b11011011;
		20'b00011110010010000110: color_data = 8'b11111111;
		20'b00011110010010000111: color_data = 8'b11111111;
		20'b00011110010010001000: color_data = 8'b11111111;
		20'b00011110010010001001: color_data = 8'b11111111;
		20'b00011110010010001010: color_data = 8'b11111111;
		20'b00011110010010001011: color_data = 8'b11111111;
		20'b00011110010010001100: color_data = 8'b11111111;
		20'b00011110010010001101: color_data = 8'b11111111;
		20'b00011110010010001110: color_data = 8'b11111111;
		20'b00011110010010011000: color_data = 8'b11011011;
		20'b00011110010010011001: color_data = 8'b11111111;
		20'b00011110010010011010: color_data = 8'b11111111;
		20'b00011110010010011011: color_data = 8'b11111111;
		20'b00011110010010011100: color_data = 8'b11111111;
		20'b00011110010010011101: color_data = 8'b11111111;
		20'b00011110010010011110: color_data = 8'b11111111;
		20'b00011110010010011111: color_data = 8'b11111111;
		20'b00011110010010100000: color_data = 8'b11111111;
		20'b00011110010010100001: color_data = 8'b11111111;
		20'b00011110010010100010: color_data = 8'b11111111;
		20'b00011110010010100011: color_data = 8'b11111111;
		20'b00011110010010100100: color_data = 8'b11111111;
		20'b00011110010010100101: color_data = 8'b11111111;
		20'b00011110010010100110: color_data = 8'b11111111;
		20'b00011110010010100111: color_data = 8'b11111111;
		20'b00011110010010101000: color_data = 8'b11111111;
		20'b00011110010010101001: color_data = 8'b11111111;
		20'b00011110010010101010: color_data = 8'b11111111;
		20'b00011110010010101011: color_data = 8'b11111111;
		20'b00011110010010101100: color_data = 8'b11111111;
		20'b00011110010010101101: color_data = 8'b11111111;
		20'b00011110010010101110: color_data = 8'b11111111;
		20'b00011110010010101111: color_data = 8'b11111111;
		20'b00011110010010110000: color_data = 8'b11111111;
		20'b00011110010010110001: color_data = 8'b11111111;
		20'b00011110010010110010: color_data = 8'b11111111;
		20'b00011110010010110011: color_data = 8'b11111111;
		20'b00011110010010110100: color_data = 8'b11111111;
		20'b00011110010010110101: color_data = 8'b11111111;
		20'b00011110010010110110: color_data = 8'b11111111;
		20'b00011110010010110111: color_data = 8'b11111111;
		20'b00011110010010111000: color_data = 8'b11111111;
		20'b00011110010010111001: color_data = 8'b11111111;
		20'b00011110010010111010: color_data = 8'b11111111;
		20'b00011110010010111011: color_data = 8'b11111111;
		20'b00011110010010111100: color_data = 8'b11111111;
		20'b00011110010010111101: color_data = 8'b11111111;
		20'b00011110010010111110: color_data = 8'b11011011;

		20'b00011110100000001001: color_data = 8'b11011011;
		20'b00011110100000001010: color_data = 8'b11111111;
		20'b00011110100000001011: color_data = 8'b11111111;
		20'b00011110100000001100: color_data = 8'b11111111;
		20'b00011110100000001101: color_data = 8'b11111111;
		20'b00011110100000001110: color_data = 8'b11111111;
		20'b00011110100000001111: color_data = 8'b11111111;
		20'b00011110100000010000: color_data = 8'b11111111;
		20'b00011110100000010001: color_data = 8'b11111111;
		20'b00011110100000010010: color_data = 8'b11111111;
		20'b00011110100000010011: color_data = 8'b10010010;
		20'b00011110100000111001: color_data = 8'b11111111;
		20'b00011110100000111010: color_data = 8'b11111111;
		20'b00011110100000111011: color_data = 8'b11111111;
		20'b00011110100000111100: color_data = 8'b11111111;
		20'b00011110100000111101: color_data = 8'b11111111;
		20'b00011110100000111110: color_data = 8'b11111111;
		20'b00011110100000111111: color_data = 8'b11111111;
		20'b00011110100001000000: color_data = 8'b11111111;
		20'b00011110100001000001: color_data = 8'b11111111;
		20'b00011110100001000010: color_data = 8'b11111111;
		20'b00011110100001000011: color_data = 8'b11111111;
		20'b00011110100001000100: color_data = 8'b11111111;
		20'b00011110100001000101: color_data = 8'b11111111;
		20'b00011110100001000110: color_data = 8'b11111111;
		20'b00011110100001000111: color_data = 8'b11111111;
		20'b00011110100001001000: color_data = 8'b11111111;
		20'b00011110100001001001: color_data = 8'b11111111;
		20'b00011110100001001010: color_data = 8'b11111111;
		20'b00011110100001001011: color_data = 8'b11111111;
		20'b00011110100001001100: color_data = 8'b11111111;
		20'b00011110100001001101: color_data = 8'b11111111;
		20'b00011110100001001110: color_data = 8'b11111111;
		20'b00011110100001001111: color_data = 8'b11111111;
		20'b00011110100001010000: color_data = 8'b11111111;
		20'b00011110100001010001: color_data = 8'b11111111;
		20'b00011110100001010010: color_data = 8'b11111111;
		20'b00011110100001010011: color_data = 8'b11111111;
		20'b00011110100001010100: color_data = 8'b11111111;
		20'b00011110100001010101: color_data = 8'b11111111;
		20'b00011110100001010110: color_data = 8'b11111111;
		20'b00011110100001010111: color_data = 8'b11111111;
		20'b00011110100001011000: color_data = 8'b11111111;
		20'b00011110100001011001: color_data = 8'b11111111;
		20'b00011110100001011010: color_data = 8'b11111111;
		20'b00011110100001011011: color_data = 8'b11111111;
		20'b00011110100001011100: color_data = 8'b11111111;
		20'b00011110100001011101: color_data = 8'b11111111;
		20'b00011110100001011110: color_data = 8'b11111111;
		20'b00011110100001011111: color_data = 8'b10010010;
		20'b00011110100001101000: color_data = 8'b10010010;
		20'b00011110100001101001: color_data = 8'b11111111;
		20'b00011110100001101010: color_data = 8'b11111111;
		20'b00011110100001101011: color_data = 8'b11111111;
		20'b00011110100001101100: color_data = 8'b11111111;
		20'b00011110100001101101: color_data = 8'b11111111;
		20'b00011110100001101110: color_data = 8'b11111111;
		20'b00011110100001101111: color_data = 8'b11111111;
		20'b00011110100001110000: color_data = 8'b11111111;
		20'b00011110100001110001: color_data = 8'b11111111;
		20'b00011110100001110010: color_data = 8'b10010010;
		20'b00011110100010000101: color_data = 8'b11011011;
		20'b00011110100010000110: color_data = 8'b11111111;
		20'b00011110100010000111: color_data = 8'b11111111;
		20'b00011110100010001000: color_data = 8'b11111111;
		20'b00011110100010001001: color_data = 8'b11111111;
		20'b00011110100010001010: color_data = 8'b11111111;
		20'b00011110100010001011: color_data = 8'b11111111;
		20'b00011110100010001100: color_data = 8'b11111111;
		20'b00011110100010001101: color_data = 8'b11111111;
		20'b00011110100010001110: color_data = 8'b11111111;
		20'b00011110100010011000: color_data = 8'b11011011;
		20'b00011110100010011001: color_data = 8'b11111111;
		20'b00011110100010011010: color_data = 8'b11111111;
		20'b00011110100010011011: color_data = 8'b11111111;
		20'b00011110100010011100: color_data = 8'b11111111;
		20'b00011110100010011101: color_data = 8'b11111111;
		20'b00011110100010011110: color_data = 8'b11111111;
		20'b00011110100010011111: color_data = 8'b11111111;
		20'b00011110100010100000: color_data = 8'b11111111;
		20'b00011110100010100001: color_data = 8'b11111111;
		20'b00011110100010100010: color_data = 8'b11111111;
		20'b00011110100010100011: color_data = 8'b11111111;
		20'b00011110100010100100: color_data = 8'b11111111;
		20'b00011110100010100101: color_data = 8'b11111111;
		20'b00011110100010100110: color_data = 8'b11111111;
		20'b00011110100010100111: color_data = 8'b11111111;
		20'b00011110100010101000: color_data = 8'b11111111;
		20'b00011110100010101001: color_data = 8'b11111111;
		20'b00011110100010101010: color_data = 8'b11111111;
		20'b00011110100010101011: color_data = 8'b11111111;
		20'b00011110100010101100: color_data = 8'b11111111;
		20'b00011110100010101101: color_data = 8'b11111111;
		20'b00011110100010101110: color_data = 8'b11111111;
		20'b00011110100010101111: color_data = 8'b11111111;
		20'b00011110100010110000: color_data = 8'b11111111;
		20'b00011110100010110001: color_data = 8'b11111111;
		20'b00011110100010110010: color_data = 8'b11111111;
		20'b00011110100010110011: color_data = 8'b11111111;
		20'b00011110100010110100: color_data = 8'b11111111;
		20'b00011110100010110101: color_data = 8'b11111111;
		20'b00011110100010110110: color_data = 8'b11111111;
		20'b00011110100010110111: color_data = 8'b11111111;
		20'b00011110100010111000: color_data = 8'b11111111;
		20'b00011110100010111001: color_data = 8'b11111111;
		20'b00011110100010111010: color_data = 8'b11111111;
		20'b00011110100010111011: color_data = 8'b11111111;
		20'b00011110100010111100: color_data = 8'b11111111;
		20'b00011110100010111101: color_data = 8'b11111111;
		20'b00011110100010111110: color_data = 8'b11011011;

		20'b00011110110000001001: color_data = 8'b11011011;
		20'b00011110110000001010: color_data = 8'b11011011;
		20'b00011110110000001011: color_data = 8'b11011011;
		20'b00011110110000001100: color_data = 8'b11011011;
		20'b00011110110000001101: color_data = 8'b11011011;
		20'b00011110110000001110: color_data = 8'b11011011;
		20'b00011110110000001111: color_data = 8'b11011011;
		20'b00011110110000010000: color_data = 8'b11011011;
		20'b00011110110000010001: color_data = 8'b11011011;
		20'b00011110110000010010: color_data = 8'b11011011;
		20'b00011110110000010011: color_data = 8'b10010010;
		20'b00011110110000111001: color_data = 8'b11011011;
		20'b00011110110000111010: color_data = 8'b11011011;
		20'b00011110110000111011: color_data = 8'b11011011;
		20'b00011110110000111100: color_data = 8'b11011011;
		20'b00011110110000111101: color_data = 8'b11011011;
		20'b00011110110000111110: color_data = 8'b11011011;
		20'b00011110110000111111: color_data = 8'b11011011;
		20'b00011110110001000000: color_data = 8'b11011011;
		20'b00011110110001000001: color_data = 8'b11011011;
		20'b00011110110001000010: color_data = 8'b11011011;
		20'b00011110110001000011: color_data = 8'b11011011;
		20'b00011110110001000100: color_data = 8'b11011011;
		20'b00011110110001000101: color_data = 8'b11011011;
		20'b00011110110001000110: color_data = 8'b11011011;
		20'b00011110110001000111: color_data = 8'b11011011;
		20'b00011110110001001000: color_data = 8'b11011011;
		20'b00011110110001001001: color_data = 8'b11011011;
		20'b00011110110001001010: color_data = 8'b11011011;
		20'b00011110110001001011: color_data = 8'b11011011;
		20'b00011110110001001100: color_data = 8'b11011011;
		20'b00011110110001001101: color_data = 8'b11011011;
		20'b00011110110001001110: color_data = 8'b11011011;
		20'b00011110110001001111: color_data = 8'b11011011;
		20'b00011110110001010000: color_data = 8'b11011011;
		20'b00011110110001010001: color_data = 8'b11011011;
		20'b00011110110001010010: color_data = 8'b11011011;
		20'b00011110110001010011: color_data = 8'b11011011;
		20'b00011110110001010100: color_data = 8'b11011011;
		20'b00011110110001010101: color_data = 8'b11011011;
		20'b00011110110001010110: color_data = 8'b11011011;
		20'b00011110110001010111: color_data = 8'b11011011;
		20'b00011110110001011000: color_data = 8'b11011011;
		20'b00011110110001011001: color_data = 8'b11011011;
		20'b00011110110001011010: color_data = 8'b11011011;
		20'b00011110110001011011: color_data = 8'b11011011;
		20'b00011110110001011100: color_data = 8'b11011011;
		20'b00011110110001011101: color_data = 8'b11011011;
		20'b00011110110001011110: color_data = 8'b11011011;
		20'b00011110110001011111: color_data = 8'b10010010;
		20'b00011110110001101000: color_data = 8'b10010010;
		20'b00011110110001101001: color_data = 8'b11011011;
		20'b00011110110001101010: color_data = 8'b11011011;
		20'b00011110110001101011: color_data = 8'b11011011;
		20'b00011110110001101100: color_data = 8'b11011011;
		20'b00011110110001101101: color_data = 8'b11011011;
		20'b00011110110001101110: color_data = 8'b11011011;
		20'b00011110110001101111: color_data = 8'b11011011;
		20'b00011110110001110000: color_data = 8'b11011011;
		20'b00011110110001110001: color_data = 8'b11011011;
		20'b00011110110001110010: color_data = 8'b10010010;
		20'b00011110110010000101: color_data = 8'b11011011;
		20'b00011110110010000110: color_data = 8'b11011011;
		20'b00011110110010000111: color_data = 8'b11011011;
		20'b00011110110010001000: color_data = 8'b11011011;
		20'b00011110110010001001: color_data = 8'b11011011;
		20'b00011110110010001010: color_data = 8'b11011011;
		20'b00011110110010001011: color_data = 8'b11011011;
		20'b00011110110010001100: color_data = 8'b11011011;
		20'b00011110110010001101: color_data = 8'b11011011;
		20'b00011110110010001110: color_data = 8'b11011011;
		20'b00011110110010011000: color_data = 8'b11011011;
		20'b00011110110010011001: color_data = 8'b11011011;
		20'b00011110110010011010: color_data = 8'b11011011;
		20'b00011110110010011011: color_data = 8'b11011011;
		20'b00011110110010011100: color_data = 8'b11011011;
		20'b00011110110010011101: color_data = 8'b11011011;
		20'b00011110110010011110: color_data = 8'b11011011;
		20'b00011110110010011111: color_data = 8'b11011011;
		20'b00011110110010100000: color_data = 8'b11011011;
		20'b00011110110010100001: color_data = 8'b11011011;
		20'b00011110110010100010: color_data = 8'b11011011;
		20'b00011110110010100011: color_data = 8'b11011011;
		20'b00011110110010100100: color_data = 8'b11011011;
		20'b00011110110010100101: color_data = 8'b11011011;
		20'b00011110110010100110: color_data = 8'b11011011;
		20'b00011110110010100111: color_data = 8'b11011011;
		20'b00011110110010101000: color_data = 8'b11011011;
		20'b00011110110010101001: color_data = 8'b11011011;
		20'b00011110110010101010: color_data = 8'b11011011;
		20'b00011110110010101011: color_data = 8'b11011011;
		20'b00011110110010101100: color_data = 8'b11011011;
		20'b00011110110010101101: color_data = 8'b11011011;
		20'b00011110110010101110: color_data = 8'b11011011;
		20'b00011110110010101111: color_data = 8'b11011011;
		20'b00011110110010110000: color_data = 8'b11011011;
		20'b00011110110010110001: color_data = 8'b11011011;
		20'b00011110110010110010: color_data = 8'b11011011;
		20'b00011110110010110011: color_data = 8'b11011011;
		20'b00011110110010110100: color_data = 8'b11011011;
		20'b00011110110010110101: color_data = 8'b11011011;
		20'b00011110110010110110: color_data = 8'b11011011;
		20'b00011110110010110111: color_data = 8'b11011011;
		20'b00011110110010111000: color_data = 8'b11011011;
		20'b00011110110010111001: color_data = 8'b11011011;
		20'b00011110110010111010: color_data = 8'b11011011;
		20'b00011110110010111011: color_data = 8'b11011011;
		20'b00011110110010111100: color_data = 8'b11011011;
		20'b00011110110010111101: color_data = 8'b11011011;
		20'b00011110110010111110: color_data = 8'b11011011;

		20'b00100111010010010011: color_data = 8'b10010010;
		20'b00100111010010010100: color_data = 8'b11111111;
		20'b00100111010010010101: color_data = 8'b11111111;
		20'b00100111010010010110: color_data = 8'b11111111;
		20'b00100111010010010111: color_data = 8'b11111111;
		20'b00100111010010011000: color_data = 8'b11111111;
		20'b00100111010010011001: color_data = 8'b11111111;
		20'b00100111010010011010: color_data = 8'b11111111;
		20'b00100111010010011011: color_data = 8'b11111111;
		20'b00100111010010011100: color_data = 8'b11111111;

		20'b00100111100010010011: color_data = 8'b10010010;
		20'b00100111100010010100: color_data = 8'b11111111;
		20'b00100111100010010101: color_data = 8'b11111111;
		20'b00100111100010010110: color_data = 8'b11111111;
		20'b00100111100010010111: color_data = 8'b11111111;
		20'b00100111100010011000: color_data = 8'b11111111;
		20'b00100111100010011001: color_data = 8'b11111111;
		20'b00100111100010011010: color_data = 8'b11111111;
		20'b00100111100010011011: color_data = 8'b11111111;
		20'b00100111100010011100: color_data = 8'b11111111;

		20'b00100111110010010011: color_data = 8'b10010010;
		20'b00100111110010010100: color_data = 8'b11111111;
		20'b00100111110010010101: color_data = 8'b11111111;
		20'b00100111110010010110: color_data = 8'b11111111;
		20'b00100111110010010111: color_data = 8'b11111111;
		20'b00100111110010011000: color_data = 8'b11111111;
		20'b00100111110010011001: color_data = 8'b11111111;
		20'b00100111110010011010: color_data = 8'b11111111;
		20'b00100111110010011011: color_data = 8'b11111111;
		20'b00100111110010011100: color_data = 8'b11111111;

		20'b00101000000010010011: color_data = 8'b10010010;
		20'b00101000000010010100: color_data = 8'b11111111;
		20'b00101000000010010101: color_data = 8'b11111111;
		20'b00101000000010010110: color_data = 8'b11111111;
		20'b00101000000010010111: color_data = 8'b11111111;
		20'b00101000000010011000: color_data = 8'b11111111;
		20'b00101000000010011001: color_data = 8'b11111111;
		20'b00101000000010011010: color_data = 8'b11111111;
		20'b00101000000010011011: color_data = 8'b11111111;
		20'b00101000000010011100: color_data = 8'b11111111;

		20'b00101000010010010011: color_data = 8'b10010010;
		20'b00101000010010010100: color_data = 8'b11111111;
		20'b00101000010010010101: color_data = 8'b11111111;
		20'b00101000010010010110: color_data = 8'b11111111;
		20'b00101000010010010111: color_data = 8'b11111111;
		20'b00101000010010011000: color_data = 8'b11111111;
		20'b00101000010010011001: color_data = 8'b11111111;
		20'b00101000010010011010: color_data = 8'b11111111;
		20'b00101000010010011011: color_data = 8'b11111111;
		20'b00101000010010011100: color_data = 8'b11111111;

		20'b00101000100010010011: color_data = 8'b10010010;
		20'b00101000100010010100: color_data = 8'b11111111;
		20'b00101000100010010101: color_data = 8'b11111111;
		20'b00101000100010010110: color_data = 8'b11111111;
		20'b00101000100010010111: color_data = 8'b11111111;
		20'b00101000100010011000: color_data = 8'b11111111;
		20'b00101000100010011001: color_data = 8'b11111111;
		20'b00101000100010011010: color_data = 8'b11111111;
		20'b00101000100010011011: color_data = 8'b11111111;
		20'b00101000100010011100: color_data = 8'b11111111;

		20'b00101000110010010011: color_data = 8'b10010010;
		20'b00101000110010010100: color_data = 8'b11111111;
		20'b00101000110010010101: color_data = 8'b11111111;
		20'b00101000110010010110: color_data = 8'b11111111;
		20'b00101000110010010111: color_data = 8'b11111111;
		20'b00101000110010011000: color_data = 8'b11111111;
		20'b00101000110010011001: color_data = 8'b11111111;
		20'b00101000110010011010: color_data = 8'b11111111;
		20'b00101000110010011011: color_data = 8'b11111111;
		20'b00101000110010011100: color_data = 8'b11111111;

		20'b00101001000010010011: color_data = 8'b10010010;
		20'b00101001000010010100: color_data = 8'b11111111;
		20'b00101001000010010101: color_data = 8'b11111111;
		20'b00101001000010010110: color_data = 8'b11111111;
		20'b00101001000010010111: color_data = 8'b11111111;
		20'b00101001000010011000: color_data = 8'b11111111;
		20'b00101001000010011001: color_data = 8'b11111111;
		20'b00101001000010011010: color_data = 8'b11111111;
		20'b00101001000010011011: color_data = 8'b11111111;
		20'b00101001000010011100: color_data = 8'b11111111;

		20'b00101001010010010011: color_data = 8'b10010010;
		20'b00101001010010010100: color_data = 8'b11111111;
		20'b00101001010010010101: color_data = 8'b11111111;
		20'b00101001010010010110: color_data = 8'b11111111;
		20'b00101001010010010111: color_data = 8'b11111111;
		20'b00101001010010011000: color_data = 8'b11111111;
		20'b00101001010010011001: color_data = 8'b11111111;
		20'b00101001010010011010: color_data = 8'b11111111;
		20'b00101001010010011011: color_data = 8'b11111111;
		20'b00101001010010011100: color_data = 8'b11111111;

		20'b00101001100010010011: color_data = 8'b10010010;
		20'b00101001100010010100: color_data = 8'b11011011;
		20'b00101001100010010101: color_data = 8'b11011011;
		20'b00101001100010010110: color_data = 8'b11011011;
		20'b00101001100010010111: color_data = 8'b11011011;
		20'b00101001100010011000: color_data = 8'b11011011;
		20'b00101001100010011001: color_data = 8'b11011011;
		20'b00101001100010011010: color_data = 8'b11011011;
		20'b00101001100010011011: color_data = 8'b11011011;
		20'b00101001100010011100: color_data = 8'b11011011;

		20'b00101101000001111100: color_data = 8'b10010010;
		20'b00101101000001111101: color_data = 8'b10010010;
		20'b00101101000001111110: color_data = 8'b10010010;
		20'b00101101000001111111: color_data = 8'b10010010;
		20'b00101101000010000000: color_data = 8'b10010010;
		20'b00101101000010000001: color_data = 8'b10010010;
		20'b00101101000010000010: color_data = 8'b10010010;
		20'b00101101000010000011: color_data = 8'b10010010;
		20'b00101101000010000100: color_data = 8'b10010010;
		20'b00101101000010000101: color_data = 8'b10010010;
		20'b00101101000010000110: color_data = 8'b10010010;
		20'b00101101000010000111: color_data = 8'b10010010;
		20'b00101101000010001000: color_data = 8'b10010010;
		20'b00101101000010001001: color_data = 8'b10010010;
		20'b00101101000010001010: color_data = 8'b10010010;
		20'b00101101000010001011: color_data = 8'b10010010;
		20'b00101101000010001100: color_data = 8'b10010010;
		20'b00101101000010001101: color_data = 8'b10010010;
		20'b00101101000010001110: color_data = 8'b10010010;
		20'b00101101000010001111: color_data = 8'b10010010;
		20'b00101101000010010000: color_data = 8'b10010010;
		20'b00101101000010010001: color_data = 8'b10010010;
		20'b00101101000010010010: color_data = 8'b10010010;
		20'b00101101000010010011: color_data = 8'b10010010;
		20'b00101101000010010100: color_data = 8'b10010010;
		20'b00101101000010010101: color_data = 8'b10010010;
		20'b00101101000010010110: color_data = 8'b10010010;
		20'b00101101000010010111: color_data = 8'b10010010;
		20'b00101101000010011000: color_data = 8'b10010010;
		20'b00101101000010011001: color_data = 8'b10010010;
		20'b00101101000010011010: color_data = 8'b10010010;
		20'b00101101000010011011: color_data = 8'b10010010;
		20'b00101101000010011100: color_data = 8'b10010010;
		20'b00101101000010011101: color_data = 8'b10010010;
		20'b00101101000010011110: color_data = 8'b10010010;
		20'b00101101000010011111: color_data = 8'b10010010;
		20'b00101101000010100000: color_data = 8'b10010010;
		20'b00101101000010100001: color_data = 8'b10010010;
		20'b00101101000010100010: color_data = 8'b10010010;
		20'b00101101000010100011: color_data = 8'b10010010;
		20'b00101101000010100100: color_data = 8'b10010010;
		20'b00101101000010100101: color_data = 8'b10010010;
		20'b00101101000010100110: color_data = 8'b10010010;
		20'b00101101000010100111: color_data = 8'b10010010;
		20'b00101101000010101000: color_data = 8'b10010010;
		20'b00101101000010101001: color_data = 8'b10010010;
		20'b00101101000010101010: color_data = 8'b10010010;
		20'b00101101000010101011: color_data = 8'b10010010;

		20'b00101101010001111011: color_data = 8'b10010010;
		20'b00101101010001111100: color_data = 8'b11011011;
		20'b00101101010001111101: color_data = 8'b11111111;
		20'b00101101010001111110: color_data = 8'b11111111;
		20'b00101101010001111111: color_data = 8'b11111111;
		20'b00101101010010000000: color_data = 8'b11111111;
		20'b00101101010010000001: color_data = 8'b11111111;
		20'b00101101010010000010: color_data = 8'b11111111;
		20'b00101101010010000011: color_data = 8'b11111111;
		20'b00101101010010000100: color_data = 8'b11111111;
		20'b00101101010010000101: color_data = 8'b11111111;
		20'b00101101010010000110: color_data = 8'b11111111;
		20'b00101101010010000111: color_data = 8'b11111111;
		20'b00101101010010001000: color_data = 8'b11111111;
		20'b00101101010010001001: color_data = 8'b11111111;
		20'b00101101010010001010: color_data = 8'b11111111;
		20'b00101101010010001011: color_data = 8'b11111111;
		20'b00101101010010001100: color_data = 8'b11111111;
		20'b00101101010010001101: color_data = 8'b11111111;
		20'b00101101010010001110: color_data = 8'b11111111;
		20'b00101101010010001111: color_data = 8'b11111111;
		20'b00101101010010010000: color_data = 8'b11111111;
		20'b00101101010010010001: color_data = 8'b11111111;
		20'b00101101010010010010: color_data = 8'b11111111;
		20'b00101101010010010011: color_data = 8'b11111111;
		20'b00101101010010010100: color_data = 8'b11111111;
		20'b00101101010010010101: color_data = 8'b11111111;
		20'b00101101010010010110: color_data = 8'b11111111;
		20'b00101101010010010111: color_data = 8'b11111111;
		20'b00101101010010011000: color_data = 8'b11111111;
		20'b00101101010010011001: color_data = 8'b11111111;
		20'b00101101010010011010: color_data = 8'b11111111;
		20'b00101101010010011011: color_data = 8'b11111111;
		20'b00101101010010011100: color_data = 8'b11111111;
		20'b00101101010010011101: color_data = 8'b11111111;
		20'b00101101010010011110: color_data = 8'b11111111;
		20'b00101101010010011111: color_data = 8'b11111111;
		20'b00101101010010100000: color_data = 8'b11111111;
		20'b00101101010010100001: color_data = 8'b11111111;
		20'b00101101010010100010: color_data = 8'b11111111;
		20'b00101101010010100011: color_data = 8'b11111111;
		20'b00101101010010100100: color_data = 8'b11111111;
		20'b00101101010010100101: color_data = 8'b11111111;
		20'b00101101010010100110: color_data = 8'b11111111;
		20'b00101101010010100111: color_data = 8'b11111111;
		20'b00101101010010101000: color_data = 8'b11111111;
		20'b00101101010010101001: color_data = 8'b11111111;
		20'b00101101010010101010: color_data = 8'b11111111;
		20'b00101101010010101011: color_data = 8'b10010010;

		20'b00101101100001111011: color_data = 8'b10010010;
		20'b00101101100001111100: color_data = 8'b11111111;
		20'b00101101100001111101: color_data = 8'b11111111;
		20'b00101101100001111110: color_data = 8'b11111111;
		20'b00101101100001111111: color_data = 8'b11111111;
		20'b00101101100010000000: color_data = 8'b11111111;
		20'b00101101100010000001: color_data = 8'b11111111;
		20'b00101101100010000010: color_data = 8'b11111111;
		20'b00101101100010000011: color_data = 8'b11111111;
		20'b00101101100010000100: color_data = 8'b11111111;
		20'b00101101100010000101: color_data = 8'b11111111;
		20'b00101101100010000110: color_data = 8'b11111111;
		20'b00101101100010000111: color_data = 8'b11111111;
		20'b00101101100010001000: color_data = 8'b11111111;
		20'b00101101100010001001: color_data = 8'b11111111;
		20'b00101101100010001010: color_data = 8'b11111111;
		20'b00101101100010001011: color_data = 8'b11111111;
		20'b00101101100010001100: color_data = 8'b11111111;
		20'b00101101100010001101: color_data = 8'b11111111;
		20'b00101101100010001110: color_data = 8'b11111111;
		20'b00101101100010001111: color_data = 8'b11111111;
		20'b00101101100010010000: color_data = 8'b11111111;
		20'b00101101100010010001: color_data = 8'b11111111;
		20'b00101101100010010010: color_data = 8'b11111111;
		20'b00101101100010010011: color_data = 8'b11111111;
		20'b00101101100010010100: color_data = 8'b11111111;
		20'b00101101100010010101: color_data = 8'b11111111;
		20'b00101101100010010110: color_data = 8'b11111111;
		20'b00101101100010010111: color_data = 8'b11111111;
		20'b00101101100010011000: color_data = 8'b11111111;
		20'b00101101100010011001: color_data = 8'b11111111;
		20'b00101101100010011010: color_data = 8'b11111111;
		20'b00101101100010011011: color_data = 8'b11111111;
		20'b00101101100010011100: color_data = 8'b11111111;
		20'b00101101100010011101: color_data = 8'b11111111;
		20'b00101101100010011110: color_data = 8'b11111111;
		20'b00101101100010011111: color_data = 8'b11111111;
		20'b00101101100010100000: color_data = 8'b11111111;
		20'b00101101100010100001: color_data = 8'b11111111;
		20'b00101101100010100010: color_data = 8'b11111111;
		20'b00101101100010100011: color_data = 8'b11111111;
		20'b00101101100010100100: color_data = 8'b11111111;
		20'b00101101100010100101: color_data = 8'b11111111;
		20'b00101101100010100110: color_data = 8'b11111111;
		20'b00101101100010100111: color_data = 8'b11111111;
		20'b00101101100010101000: color_data = 8'b11111111;
		20'b00101101100010101001: color_data = 8'b11111111;
		20'b00101101100010101010: color_data = 8'b11111111;
		20'b00101101100010101011: color_data = 8'b10010010;

		20'b00101101110001111011: color_data = 8'b10010010;
		20'b00101101110001111100: color_data = 8'b11111111;
		20'b00101101110001111101: color_data = 8'b11111111;
		20'b00101101110001111110: color_data = 8'b11111111;
		20'b00101101110001111111: color_data = 8'b11111111;
		20'b00101101110010000000: color_data = 8'b11111111;
		20'b00101101110010000001: color_data = 8'b11111111;
		20'b00101101110010000010: color_data = 8'b11111111;
		20'b00101101110010000011: color_data = 8'b11111111;
		20'b00101101110010000100: color_data = 8'b11111111;
		20'b00101101110010000101: color_data = 8'b11111111;
		20'b00101101110010000110: color_data = 8'b11111111;
		20'b00101101110010000111: color_data = 8'b11111111;
		20'b00101101110010001000: color_data = 8'b11111111;
		20'b00101101110010001001: color_data = 8'b11111111;
		20'b00101101110010001010: color_data = 8'b11111111;
		20'b00101101110010001011: color_data = 8'b11111111;
		20'b00101101110010001100: color_data = 8'b11111111;
		20'b00101101110010001101: color_data = 8'b11111111;
		20'b00101101110010001110: color_data = 8'b11111111;
		20'b00101101110010001111: color_data = 8'b11111111;
		20'b00101101110010010000: color_data = 8'b11111111;
		20'b00101101110010010001: color_data = 8'b11111111;
		20'b00101101110010010010: color_data = 8'b11111111;
		20'b00101101110010010011: color_data = 8'b11111111;
		20'b00101101110010010100: color_data = 8'b11111111;
		20'b00101101110010010101: color_data = 8'b11111111;
		20'b00101101110010010110: color_data = 8'b11111111;
		20'b00101101110010010111: color_data = 8'b11111111;
		20'b00101101110010011000: color_data = 8'b11111111;
		20'b00101101110010011001: color_data = 8'b11111111;
		20'b00101101110010011010: color_data = 8'b11111111;
		20'b00101101110010011011: color_data = 8'b11111111;
		20'b00101101110010011100: color_data = 8'b11111111;
		20'b00101101110010011101: color_data = 8'b11111111;
		20'b00101101110010011110: color_data = 8'b11111111;
		20'b00101101110010011111: color_data = 8'b11111111;
		20'b00101101110010100000: color_data = 8'b11111111;
		20'b00101101110010100001: color_data = 8'b11111111;
		20'b00101101110010100010: color_data = 8'b11111111;
		20'b00101101110010100011: color_data = 8'b11111111;
		20'b00101101110010100100: color_data = 8'b11111111;
		20'b00101101110010100101: color_data = 8'b11111111;
		20'b00101101110010100110: color_data = 8'b11111111;
		20'b00101101110010100111: color_data = 8'b11111111;
		20'b00101101110010101000: color_data = 8'b11111111;
		20'b00101101110010101001: color_data = 8'b11111111;
		20'b00101101110010101010: color_data = 8'b11111111;
		20'b00101101110010101011: color_data = 8'b10010010;

		20'b00101110000001111011: color_data = 8'b10010010;
		20'b00101110000001111100: color_data = 8'b11111111;
		20'b00101110000001111101: color_data = 8'b11111111;
		20'b00101110000001111110: color_data = 8'b11111111;
		20'b00101110000001111111: color_data = 8'b11111111;
		20'b00101110000010000000: color_data = 8'b11111111;
		20'b00101110000010000001: color_data = 8'b11111111;
		20'b00101110000010000010: color_data = 8'b11111111;
		20'b00101110000010000011: color_data = 8'b11111111;
		20'b00101110000010000100: color_data = 8'b11111111;
		20'b00101110000010000101: color_data = 8'b11111111;
		20'b00101110000010000110: color_data = 8'b11111111;
		20'b00101110000010000111: color_data = 8'b11111111;
		20'b00101110000010001000: color_data = 8'b11111111;
		20'b00101110000010001001: color_data = 8'b11111111;
		20'b00101110000010001010: color_data = 8'b11111111;
		20'b00101110000010001011: color_data = 8'b11111111;
		20'b00101110000010001100: color_data = 8'b11111111;
		20'b00101110000010001101: color_data = 8'b11111111;
		20'b00101110000010001110: color_data = 8'b11111111;
		20'b00101110000010001111: color_data = 8'b11111111;
		20'b00101110000010010000: color_data = 8'b11111111;
		20'b00101110000010010001: color_data = 8'b11111111;
		20'b00101110000010010010: color_data = 8'b11111111;
		20'b00101110000010010011: color_data = 8'b11111111;
		20'b00101110000010010100: color_data = 8'b11111111;
		20'b00101110000010010101: color_data = 8'b11111111;
		20'b00101110000010010110: color_data = 8'b11111111;
		20'b00101110000010010111: color_data = 8'b11111111;
		20'b00101110000010011000: color_data = 8'b11111111;
		20'b00101110000010011001: color_data = 8'b11111111;
		20'b00101110000010011010: color_data = 8'b11111111;
		20'b00101110000010011011: color_data = 8'b11111111;
		20'b00101110000010011100: color_data = 8'b11111111;
		20'b00101110000010011101: color_data = 8'b11111111;
		20'b00101110000010011110: color_data = 8'b11111111;
		20'b00101110000010011111: color_data = 8'b11111111;
		20'b00101110000010100000: color_data = 8'b11111111;
		20'b00101110000010100001: color_data = 8'b11111111;
		20'b00101110000010100010: color_data = 8'b11111111;
		20'b00101110000010100011: color_data = 8'b11111111;
		20'b00101110000010100100: color_data = 8'b11111111;
		20'b00101110000010100101: color_data = 8'b11111111;
		20'b00101110000010100110: color_data = 8'b11111111;
		20'b00101110000010100111: color_data = 8'b11111111;
		20'b00101110000010101000: color_data = 8'b11111111;
		20'b00101110000010101001: color_data = 8'b11111111;
		20'b00101110000010101010: color_data = 8'b11111111;
		20'b00101110000010101011: color_data = 8'b11011011;

		20'b00101110010001111011: color_data = 8'b10010010;
		20'b00101110010001111100: color_data = 8'b11111111;
		20'b00101110010001111101: color_data = 8'b11111111;
		20'b00101110010001111110: color_data = 8'b11111111;
		20'b00101110010001111111: color_data = 8'b11111111;
		20'b00101110010010000000: color_data = 8'b11111111;
		20'b00101110010010000001: color_data = 8'b11111111;
		20'b00101110010010000010: color_data = 8'b11111111;
		20'b00101110010010000011: color_data = 8'b11111111;
		20'b00101110010010000100: color_data = 8'b11111111;
		20'b00101110010010000101: color_data = 8'b11111111;
		20'b00101110010010000110: color_data = 8'b11111111;
		20'b00101110010010000111: color_data = 8'b11111111;
		20'b00101110010010001000: color_data = 8'b11111111;
		20'b00101110010010001001: color_data = 8'b11111111;
		20'b00101110010010001010: color_data = 8'b11111111;
		20'b00101110010010001011: color_data = 8'b11111111;
		20'b00101110010010001100: color_data = 8'b11111111;
		20'b00101110010010001101: color_data = 8'b11111111;
		20'b00101110010010001110: color_data = 8'b11111111;
		20'b00101110010010001111: color_data = 8'b11111111;
		20'b00101110010010010000: color_data = 8'b11111111;
		20'b00101110010010010001: color_data = 8'b11111111;
		20'b00101110010010010010: color_data = 8'b11111111;
		20'b00101110010010010011: color_data = 8'b11111111;
		20'b00101110010010010100: color_data = 8'b11111111;
		20'b00101110010010010101: color_data = 8'b11111111;
		20'b00101110010010010110: color_data = 8'b11111111;
		20'b00101110010010010111: color_data = 8'b11111111;
		20'b00101110010010011000: color_data = 8'b11111111;
		20'b00101110010010011001: color_data = 8'b11111111;
		20'b00101110010010011010: color_data = 8'b11111111;
		20'b00101110010010011011: color_data = 8'b11111111;
		20'b00101110010010011100: color_data = 8'b11111111;
		20'b00101110010010011101: color_data = 8'b11111111;
		20'b00101110010010011110: color_data = 8'b11111111;
		20'b00101110010010011111: color_data = 8'b11111111;
		20'b00101110010010100000: color_data = 8'b11111111;
		20'b00101110010010100001: color_data = 8'b11111111;
		20'b00101110010010100010: color_data = 8'b11111111;
		20'b00101110010010100011: color_data = 8'b11111111;
		20'b00101110010010100100: color_data = 8'b11111111;
		20'b00101110010010100101: color_data = 8'b11111111;
		20'b00101110010010100110: color_data = 8'b11111111;
		20'b00101110010010100111: color_data = 8'b11111111;
		20'b00101110010010101000: color_data = 8'b11111111;
		20'b00101110010010101001: color_data = 8'b11111111;
		20'b00101110010010101010: color_data = 8'b11111111;
		20'b00101110010010101011: color_data = 8'b10010010;

		20'b00101110100001111011: color_data = 8'b10010010;
		20'b00101110100001111100: color_data = 8'b11111111;
		20'b00101110100001111101: color_data = 8'b11111111;
		20'b00101110100001111110: color_data = 8'b11111111;
		20'b00101110100001111111: color_data = 8'b11111111;
		20'b00101110100010000000: color_data = 8'b11111111;
		20'b00101110100010000001: color_data = 8'b11111111;
		20'b00101110100010000010: color_data = 8'b11111111;
		20'b00101110100010000011: color_data = 8'b11111111;
		20'b00101110100010000100: color_data = 8'b11111111;
		20'b00101110100010000101: color_data = 8'b11111111;
		20'b00101110100010000110: color_data = 8'b11111111;
		20'b00101110100010000111: color_data = 8'b11111111;
		20'b00101110100010001000: color_data = 8'b11111111;
		20'b00101110100010001001: color_data = 8'b11111111;
		20'b00101110100010001010: color_data = 8'b11111111;
		20'b00101110100010001011: color_data = 8'b11111111;
		20'b00101110100010001100: color_data = 8'b11111111;
		20'b00101110100010001101: color_data = 8'b11111111;
		20'b00101110100010001110: color_data = 8'b11111111;
		20'b00101110100010001111: color_data = 8'b11111111;
		20'b00101110100010010000: color_data = 8'b11111111;
		20'b00101110100010010001: color_data = 8'b11111111;
		20'b00101110100010010010: color_data = 8'b11111111;
		20'b00101110100010010011: color_data = 8'b11111111;
		20'b00101110100010010100: color_data = 8'b11111111;
		20'b00101110100010010101: color_data = 8'b11111111;
		20'b00101110100010010110: color_data = 8'b11111111;
		20'b00101110100010010111: color_data = 8'b11111111;
		20'b00101110100010011000: color_data = 8'b11111111;
		20'b00101110100010011001: color_data = 8'b11111111;
		20'b00101110100010011010: color_data = 8'b11111111;
		20'b00101110100010011011: color_data = 8'b11111111;
		20'b00101110100010011100: color_data = 8'b11111111;
		20'b00101110100010011101: color_data = 8'b11111111;
		20'b00101110100010011110: color_data = 8'b11111111;
		20'b00101110100010011111: color_data = 8'b11111111;
		20'b00101110100010100000: color_data = 8'b11111111;
		20'b00101110100010100001: color_data = 8'b11111111;
		20'b00101110100010100010: color_data = 8'b11111111;
		20'b00101110100010100011: color_data = 8'b11111111;
		20'b00101110100010100100: color_data = 8'b11111111;
		20'b00101110100010100101: color_data = 8'b11111111;
		20'b00101110100010100110: color_data = 8'b11111111;
		20'b00101110100010100111: color_data = 8'b11111111;
		20'b00101110100010101000: color_data = 8'b11111111;
		20'b00101110100010101001: color_data = 8'b11111111;
		20'b00101110100010101010: color_data = 8'b11111111;
		20'b00101110100010101011: color_data = 8'b11011011;

		20'b00101110110001111011: color_data = 8'b10010010;
		20'b00101110110001111100: color_data = 8'b11111111;
		20'b00101110110001111101: color_data = 8'b11111111;
		20'b00101110110001111110: color_data = 8'b11111111;
		20'b00101110110001111111: color_data = 8'b11111111;
		20'b00101110110010000000: color_data = 8'b11111111;
		20'b00101110110010000001: color_data = 8'b11111111;
		20'b00101110110010000010: color_data = 8'b11111111;
		20'b00101110110010000011: color_data = 8'b11111111;
		20'b00101110110010000100: color_data = 8'b11111111;
		20'b00101110110010000101: color_data = 8'b11111111;
		20'b00101110110010000110: color_data = 8'b11111111;
		20'b00101110110010000111: color_data = 8'b11111111;
		20'b00101110110010001000: color_data = 8'b11111111;
		20'b00101110110010001001: color_data = 8'b11111111;
		20'b00101110110010001010: color_data = 8'b11111111;
		20'b00101110110010001011: color_data = 8'b11111111;
		20'b00101110110010001100: color_data = 8'b11111111;
		20'b00101110110010001101: color_data = 8'b11111111;
		20'b00101110110010001110: color_data = 8'b11111111;
		20'b00101110110010001111: color_data = 8'b11111111;
		20'b00101110110010010000: color_data = 8'b11111111;
		20'b00101110110010010001: color_data = 8'b11111111;
		20'b00101110110010010010: color_data = 8'b11111111;
		20'b00101110110010010011: color_data = 8'b11111111;
		20'b00101110110010010100: color_data = 8'b11111111;
		20'b00101110110010010101: color_data = 8'b11111111;
		20'b00101110110010010110: color_data = 8'b11111111;
		20'b00101110110010010111: color_data = 8'b11111111;
		20'b00101110110010011000: color_data = 8'b11111111;
		20'b00101110110010011001: color_data = 8'b11111111;
		20'b00101110110010011010: color_data = 8'b11111111;
		20'b00101110110010011011: color_data = 8'b11111111;
		20'b00101110110010011100: color_data = 8'b11111111;
		20'b00101110110010011101: color_data = 8'b11111111;
		20'b00101110110010011110: color_data = 8'b11111111;
		20'b00101110110010011111: color_data = 8'b11111111;
		20'b00101110110010100000: color_data = 8'b11111111;
		20'b00101110110010100001: color_data = 8'b11111111;
		20'b00101110110010100010: color_data = 8'b11111111;
		20'b00101110110010100011: color_data = 8'b11111111;
		20'b00101110110010100100: color_data = 8'b11111111;
		20'b00101110110010100101: color_data = 8'b11111111;
		20'b00101110110010100110: color_data = 8'b11111111;
		20'b00101110110010100111: color_data = 8'b11111111;
		20'b00101110110010101000: color_data = 8'b11111111;
		20'b00101110110010101001: color_data = 8'b11111111;
		20'b00101110110010101010: color_data = 8'b11111111;
		20'b00101110110010101011: color_data = 8'b11011011;

		20'b00101111000001111011: color_data = 8'b10010010;
		20'b00101111000001111100: color_data = 8'b11111111;
		20'b00101111000001111101: color_data = 8'b11111111;
		20'b00101111000001111110: color_data = 8'b11111111;
		20'b00101111000001111111: color_data = 8'b11111111;
		20'b00101111000010000000: color_data = 8'b11111111;
		20'b00101111000010000001: color_data = 8'b11111111;
		20'b00101111000010000010: color_data = 8'b11111111;
		20'b00101111000010000011: color_data = 8'b11111111;
		20'b00101111000010000100: color_data = 8'b11111111;
		20'b00101111000010000101: color_data = 8'b11111111;
		20'b00101111000010000110: color_data = 8'b11111111;
		20'b00101111000010000111: color_data = 8'b11111111;
		20'b00101111000010001000: color_data = 8'b11111111;
		20'b00101111000010001001: color_data = 8'b11111111;
		20'b00101111000010001010: color_data = 8'b11111111;
		20'b00101111000010001011: color_data = 8'b11111111;
		20'b00101111000010001100: color_data = 8'b11111111;
		20'b00101111000010001101: color_data = 8'b11111111;
		20'b00101111000010001110: color_data = 8'b11111111;
		20'b00101111000010001111: color_data = 8'b11111111;
		20'b00101111000010010000: color_data = 8'b11111111;
		20'b00101111000010010001: color_data = 8'b11111111;
		20'b00101111000010010010: color_data = 8'b11111111;
		20'b00101111000010010011: color_data = 8'b11111111;
		20'b00101111000010010100: color_data = 8'b11111111;
		20'b00101111000010010101: color_data = 8'b11111111;
		20'b00101111000010010110: color_data = 8'b11111111;
		20'b00101111000010010111: color_data = 8'b11111111;
		20'b00101111000010011000: color_data = 8'b11111111;
		20'b00101111000010011001: color_data = 8'b11111111;
		20'b00101111000010011010: color_data = 8'b11111111;
		20'b00101111000010011011: color_data = 8'b11111111;
		20'b00101111000010011100: color_data = 8'b11111111;
		20'b00101111000010011101: color_data = 8'b11111111;
		20'b00101111000010011110: color_data = 8'b11111111;
		20'b00101111000010011111: color_data = 8'b11111111;
		20'b00101111000010100000: color_data = 8'b11111111;
		20'b00101111000010100001: color_data = 8'b11111111;
		20'b00101111000010100010: color_data = 8'b11111111;
		20'b00101111000010100011: color_data = 8'b11111111;
		20'b00101111000010100100: color_data = 8'b11111111;
		20'b00101111000010100101: color_data = 8'b11111111;
		20'b00101111000010100110: color_data = 8'b11111111;
		20'b00101111000010100111: color_data = 8'b11111111;
		20'b00101111000010101000: color_data = 8'b11111111;
		20'b00101111000010101001: color_data = 8'b11111111;
		20'b00101111000010101010: color_data = 8'b11111111;
		20'b00101111000010101011: color_data = 8'b11011011;

		20'b00101111010001111011: color_data = 8'b10010010;
		20'b00101111010001111100: color_data = 8'b11111111;
		20'b00101111010001111101: color_data = 8'b11111111;
		20'b00101111010001111110: color_data = 8'b11111111;
		20'b00101111010001111111: color_data = 8'b11111111;
		20'b00101111010010000000: color_data = 8'b11111111;
		20'b00101111010010000001: color_data = 8'b11111111;
		20'b00101111010010000010: color_data = 8'b11111111;
		20'b00101111010010000011: color_data = 8'b11111111;
		20'b00101111010010000100: color_data = 8'b11111111;
		20'b00101111010010000101: color_data = 8'b11111111;
		20'b00101111010010000110: color_data = 8'b11111111;
		20'b00101111010010000111: color_data = 8'b11111111;
		20'b00101111010010001000: color_data = 8'b11111111;
		20'b00101111010010001001: color_data = 8'b11111111;
		20'b00101111010010001010: color_data = 8'b11111111;
		20'b00101111010010001011: color_data = 8'b11111111;
		20'b00101111010010001100: color_data = 8'b11111111;
		20'b00101111010010001101: color_data = 8'b11111111;
		20'b00101111010010001110: color_data = 8'b11111111;
		20'b00101111010010001111: color_data = 8'b11111111;
		20'b00101111010010010000: color_data = 8'b11111111;
		20'b00101111010010010001: color_data = 8'b11111111;
		20'b00101111010010010010: color_data = 8'b11111111;
		20'b00101111010010010011: color_data = 8'b11111111;
		20'b00101111010010010100: color_data = 8'b11111111;
		20'b00101111010010010101: color_data = 8'b11111111;
		20'b00101111010010010110: color_data = 8'b11111111;
		20'b00101111010010010111: color_data = 8'b11111111;
		20'b00101111010010011000: color_data = 8'b11111111;
		20'b00101111010010011001: color_data = 8'b11111111;
		20'b00101111010010011010: color_data = 8'b11111111;
		20'b00101111010010011011: color_data = 8'b11111111;
		20'b00101111010010011100: color_data = 8'b11111111;
		20'b00101111010010011101: color_data = 8'b11111111;
		20'b00101111010010011110: color_data = 8'b11111111;
		20'b00101111010010011111: color_data = 8'b11111111;
		20'b00101111010010100000: color_data = 8'b11111111;
		20'b00101111010010100001: color_data = 8'b11111111;
		20'b00101111010010100010: color_data = 8'b11111111;
		20'b00101111010010100011: color_data = 8'b11111111;
		20'b00101111010010100100: color_data = 8'b11111111;
		20'b00101111010010100101: color_data = 8'b11111111;
		20'b00101111010010100110: color_data = 8'b11111111;
		20'b00101111010010100111: color_data = 8'b11111111;
		20'b00101111010010101000: color_data = 8'b11111111;
		20'b00101111010010101001: color_data = 8'b11111111;
		20'b00101111010010101010: color_data = 8'b11111111;
		20'b00101111010010101011: color_data = 8'b11011011;

		20'b00101111100001111011: color_data = 8'b10010010;
		20'b00101111100001111100: color_data = 8'b11011011;
		20'b00101111100001111101: color_data = 8'b11011011;
		20'b00101111100001111110: color_data = 8'b11011011;
		20'b00101111100001111111: color_data = 8'b11011011;
		20'b00101111100010000000: color_data = 8'b11011011;
		20'b00101111100010000001: color_data = 8'b11011011;
		20'b00101111100010000010: color_data = 8'b11011011;
		20'b00101111100010000011: color_data = 8'b11011011;
		20'b00101111100010000100: color_data = 8'b11011011;
		20'b00101111100010000101: color_data = 8'b11011011;
		20'b00101111100010000110: color_data = 8'b11011011;
		20'b00101111100010000111: color_data = 8'b11011011;
		20'b00101111100010001000: color_data = 8'b11011011;
		20'b00101111100010001001: color_data = 8'b11011011;
		20'b00101111100010001010: color_data = 8'b11011011;
		20'b00101111100010001011: color_data = 8'b11011011;
		20'b00101111100010001100: color_data = 8'b11011011;
		20'b00101111100010001101: color_data = 8'b11011011;
		20'b00101111100010001110: color_data = 8'b11011011;
		20'b00101111100010001111: color_data = 8'b11011011;
		20'b00101111100010010000: color_data = 8'b11011011;
		20'b00101111100010010001: color_data = 8'b11011011;
		20'b00101111100010010010: color_data = 8'b11011011;
		20'b00101111100010010011: color_data = 8'b11011011;
		20'b00101111100010010100: color_data = 8'b11011011;
		20'b00101111100010010101: color_data = 8'b11011011;
		20'b00101111100010010110: color_data = 8'b11011011;
		20'b00101111100010010111: color_data = 8'b11011011;
		20'b00101111100010011000: color_data = 8'b11011011;
		20'b00101111100010011001: color_data = 8'b11011011;
		20'b00101111100010011010: color_data = 8'b11011011;
		20'b00101111100010011011: color_data = 8'b11011011;
		20'b00101111100010011100: color_data = 8'b11011011;
		20'b00101111100010011101: color_data = 8'b11011011;
		20'b00101111100010011110: color_data = 8'b11011011;
		20'b00101111100010011111: color_data = 8'b11011011;
		20'b00101111100010100000: color_data = 8'b11011011;
		20'b00101111100010100001: color_data = 8'b11011011;
		20'b00101111100010100010: color_data = 8'b11011011;
		20'b00101111100010100011: color_data = 8'b11011011;
		20'b00101111100010100100: color_data = 8'b11011011;
		20'b00101111100010100101: color_data = 8'b11011011;
		20'b00101111100010100110: color_data = 8'b11011011;
		20'b00101111100010100111: color_data = 8'b11011011;
		20'b00101111100010101000: color_data = 8'b11011011;
		20'b00101111100010101001: color_data = 8'b11011011;
		20'b00101111100010101010: color_data = 8'b11011011;
		20'b00101111100010101011: color_data = 8'b10010010;

		default: color_data = 8'b00000000;
	endcase
endmodule