////////////////////////////////////////////////////////////
//
//	Names: Larry Kozlowski and Alexander Romero
// Date: 2/22/17
// CM#1125 and CM#3297
// Purpose: Pixel colors for the pong logo
////////////////////////////////////////////////////////////

module pong_logo_rom
	(
		input wire clk,
		input wire [9:0] xpos,
		input wire [9:0] ypos,
		output reg [2:0] red,
		output reg [2:0] green,
		output reg [1:0] blue
	);

	(* rom_style = "block" *)


	reg [9:0] ypos_reg;
	reg [9:0] xpos_reg;

	always @(posedge clk)
		begin
		ypos_reg <= ypos;
		xpos_reg <= xpos;
		end

	always @*
	case ({xpos_reg, ypos_reg})
		20'b00000010010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001001101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001001111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001010000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001011101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001011110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001100000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001101011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001101100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001101101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001101110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001101111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001110000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000010110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001011101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001011110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110001101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001101011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001101100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001101101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001101110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001101111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001110000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001110001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001110010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110001111011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000101000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001001010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001011101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001011110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001001101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001001111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001010000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001011101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001011110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001100000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000001110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001101000000001111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001100000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001101011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001101100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001101101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001101110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001101111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001110000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001011101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001011110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001011111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001100000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001100001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001100010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001101011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001101100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001101101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001101110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001101111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001110000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001110001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111110001001100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001001101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001001110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001001111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001010000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001010001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001010010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001011101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001011110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001011111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001100000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001100001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001100010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001101011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001101100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001101101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001101110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001101111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001110000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001110001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001110010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111110001111011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011000000000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000010000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001001100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001001101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001001110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001001111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001010000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001010001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001010010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001011101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001011110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001011111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001100000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001100001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001100010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001101011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001101100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001101101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001101110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001101111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001110000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001110001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001110010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000001111011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001011101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001011110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001011111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001100000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001100001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001100010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001101011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001101100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001101101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001101110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001101111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001110000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001110001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001110010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100100001111011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110010110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010111011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010111100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010111101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110010111110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000010110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011111100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011111110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100000000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100000100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100000110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001100000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001101011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001101100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001101101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001101110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001101111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001110000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100011010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100011100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100011110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110010011101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010011110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010011111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010100000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010100001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010100010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100101010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100101100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001001101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001001111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001010000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001011101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001011110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001100000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001101011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001101100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001101101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001101110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001101111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001110000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110100010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000010011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100111000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100111010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100111100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100111110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101000000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001011101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001011110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001100000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001101011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001101100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001101101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001101110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001101111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001110000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101000010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101000100001110010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101000100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101000100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101000110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101001000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101001010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101001100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101001110010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010000010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010010010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010100010110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100010111110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001011111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010110001100000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110010110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010110010110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010110010110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010110010110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010110010111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110010111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010110010111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110010111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110010111100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110010111101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110010111110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101011000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001101011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001101100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001101101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001101110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001101111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001110000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001110001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101000001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110110001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110110001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110110001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110110001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001011111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001001100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001001101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001001110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001001111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001010000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101111100001011111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101111100001100000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001101011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001101100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001101101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001101110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001101111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001110000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001111011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		default: begin red <= 3'b000; green <= 3'b000; blue <= 2'b00; end
	endcase
endmodule