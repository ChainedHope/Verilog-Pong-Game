module credit_menu_rom
	(
		input wire clk,
		input wire [9:0] row,
		input wire [9:0] col,
		output reg [7:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [9:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		20'b00000001100000010101: color_data = 8'b11111111;
		20'b00000001100000010110: color_data = 8'b11111111;
		20'b00000001100000010111: color_data = 8'b11111111;
		20'b00000001100000011000: color_data = 8'b11111111;
		20'b00000001100000011001: color_data = 8'b11111111;
		20'b00000001110000010011: color_data = 8'b11111111;
		20'b00000001110000010100: color_data = 8'b11111111;
		20'b00000001110000010101: color_data = 8'b11111111;
		20'b00000001110000010110: color_data = 8'b11111111;
		20'b00000001110000010111: color_data = 8'b11111111;
		20'b00000001110000011000: color_data = 8'b11111111;
		20'b00000001110000011001: color_data = 8'b11111111;
		20'b00000001110000011010: color_data = 8'b11111111;
		20'b00000010000000010011: color_data = 8'b11111111;
		20'b00000010000000010100: color_data = 8'b11111111;
		20'b00000010000000010101: color_data = 8'b11111111;
		20'b00000010000000011010: color_data = 8'b11111111;
		20'b00000010000000011011: color_data = 8'b11111111;
		20'b00000010000000011100: color_data = 8'b11111111;
		20'b00000010000000011111: color_data = 8'b11111111;
		20'b00000010000000100000: color_data = 8'b11111111;
		20'b00000010000000100001: color_data = 8'b11111111;
		20'b00000010000000100010: color_data = 8'b11111111;
		20'b00000010000000100011: color_data = 8'b11111111;
		20'b00000010000000100100: color_data = 8'b11111111;
		20'b00000010000000100101: color_data = 8'b11111111;
		20'b00000010000000101001: color_data = 8'b11111111;
		20'b00000010000000101010: color_data = 8'b11111111;
		20'b00000010000000101011: color_data = 8'b11111111;
		20'b00000010000000101100: color_data = 8'b11111111;
		20'b00000010000000101101: color_data = 8'b11111111;
		20'b00000010000000101110: color_data = 8'b11111111;
		20'b00000010000000101111: color_data = 8'b11111111;
		20'b00000010000000110000: color_data = 8'b11111111;
		20'b00000010000000110011: color_data = 8'b11111111;
		20'b00000010000000110100: color_data = 8'b11111111;
		20'b00000010000000110101: color_data = 8'b11111111;
		20'b00000010000000110110: color_data = 8'b11111111;
		20'b00000010000000110111: color_data = 8'b11111111;
		20'b00000010000000111000: color_data = 8'b11111111;
		20'b00000010000000111001: color_data = 8'b11111111;
		20'b00000010000000111110: color_data = 8'b11111111;
		20'b00000010000000111111: color_data = 8'b11111111;
		20'b00000010000001000001: color_data = 8'b11111111;
		20'b00000010000001000010: color_data = 8'b11111111;
		20'b00000010000001000011: color_data = 8'b11111111;
		20'b00000010000001000100: color_data = 8'b11111111;
		20'b00000010000001000101: color_data = 8'b11111111;
		20'b00000010000001000110: color_data = 8'b11111111;
		20'b00000010000001000111: color_data = 8'b11111111;
		20'b00000010000001001000: color_data = 8'b11111111;
		20'b00000010000001001100: color_data = 8'b11111111;
		20'b00000010000001001101: color_data = 8'b11111111;
		20'b00000010000001001110: color_data = 8'b11111111;
		20'b00000010000001001111: color_data = 8'b11111111;
		20'b00000010010000010010: color_data = 8'b11111111;
		20'b00000010010000010011: color_data = 8'b11111111;
		20'b00000010010000011011: color_data = 8'b11111111;
		20'b00000010010000011111: color_data = 8'b11111111;
		20'b00000010010000100000: color_data = 8'b11111111;
		20'b00000010010000100001: color_data = 8'b11111111;
		20'b00000010010000100010: color_data = 8'b11111111;
		20'b00000010010000100011: color_data = 8'b11111111;
		20'b00000010010000100100: color_data = 8'b11111111;
		20'b00000010010000100101: color_data = 8'b11111111;
		20'b00000010010000100110: color_data = 8'b11111111;
		20'b00000010010000101001: color_data = 8'b11111111;
		20'b00000010010000101010: color_data = 8'b11111111;
		20'b00000010010000101011: color_data = 8'b11111111;
		20'b00000010010000101100: color_data = 8'b11111111;
		20'b00000010010000101101: color_data = 8'b11111111;
		20'b00000010010000101110: color_data = 8'b11111111;
		20'b00000010010000101111: color_data = 8'b11111111;
		20'b00000010010000110000: color_data = 8'b11111111;
		20'b00000010010000110011: color_data = 8'b11111111;
		20'b00000010010000110100: color_data = 8'b11111111;
		20'b00000010010000110101: color_data = 8'b11111111;
		20'b00000010010000110110: color_data = 8'b11111111;
		20'b00000010010000110111: color_data = 8'b11111111;
		20'b00000010010000111000: color_data = 8'b11111111;
		20'b00000010010000111001: color_data = 8'b11111111;
		20'b00000010010000111010: color_data = 8'b11111111;
		20'b00000010010000111110: color_data = 8'b11111111;
		20'b00000010010000111111: color_data = 8'b11111111;
		20'b00000010010001000001: color_data = 8'b11111111;
		20'b00000010010001000010: color_data = 8'b11111111;
		20'b00000010010001000011: color_data = 8'b11111111;
		20'b00000010010001000100: color_data = 8'b11111111;
		20'b00000010010001000101: color_data = 8'b11111111;
		20'b00000010010001000110: color_data = 8'b11111111;
		20'b00000010010001000111: color_data = 8'b11111111;
		20'b00000010010001001000: color_data = 8'b11111111;
		20'b00000010010001001011: color_data = 8'b11111111;
		20'b00000010010001001100: color_data = 8'b11111111;
		20'b00000010010001001101: color_data = 8'b11111111;
		20'b00000010010001001110: color_data = 8'b11111111;
		20'b00000010010001001111: color_data = 8'b11111111;
		20'b00000010010001010000: color_data = 8'b11111111;
		20'b00000010010001010001: color_data = 8'b11111111;
		20'b00000010100000010010: color_data = 8'b11111111;
		20'b00000010100000010011: color_data = 8'b11111111;
		20'b00000010100000011111: color_data = 8'b11111111;
		20'b00000010100000100000: color_data = 8'b11111111;
		20'b00000010100000100101: color_data = 8'b11111111;
		20'b00000010100000100110: color_data = 8'b11111111;
		20'b00000010100000101001: color_data = 8'b11111111;
		20'b00000010100000101010: color_data = 8'b11111111;
		20'b00000010100000110011: color_data = 8'b11111111;
		20'b00000010100000110100: color_data = 8'b11111111;
		20'b00000010100000111001: color_data = 8'b11111111;
		20'b00000010100000111010: color_data = 8'b11111111;
		20'b00000010100000111011: color_data = 8'b11111111;
		20'b00000010100000111110: color_data = 8'b11111111;
		20'b00000010100000111111: color_data = 8'b11111111;
		20'b00000010100001000100: color_data = 8'b11111111;
		20'b00000010100001000101: color_data = 8'b11111111;
		20'b00000010100001001011: color_data = 8'b11111111;
		20'b00000010100001001100: color_data = 8'b11111111;
		20'b00000010100001010001: color_data = 8'b11111111;
		20'b00000010110000010010: color_data = 8'b11111111;
		20'b00000010110000010011: color_data = 8'b11111111;
		20'b00000010110000011111: color_data = 8'b11111111;
		20'b00000010110000100000: color_data = 8'b11111111;
		20'b00000010110000100001: color_data = 8'b11111111;
		20'b00000010110000100010: color_data = 8'b11111111;
		20'b00000010110000100011: color_data = 8'b11111111;
		20'b00000010110000100100: color_data = 8'b11111111;
		20'b00000010110000100101: color_data = 8'b11111111;
		20'b00000010110000100110: color_data = 8'b11111111;
		20'b00000010110000101001: color_data = 8'b11111111;
		20'b00000010110000101010: color_data = 8'b11111111;
		20'b00000010110000101011: color_data = 8'b11111111;
		20'b00000010110000101100: color_data = 8'b11111111;
		20'b00000010110000101101: color_data = 8'b11111111;
		20'b00000010110000101110: color_data = 8'b11111111;
		20'b00000010110000110011: color_data = 8'b11111111;
		20'b00000010110000110100: color_data = 8'b11111111;
		20'b00000010110000111010: color_data = 8'b11111111;
		20'b00000010110000111011: color_data = 8'b11111111;
		20'b00000010110000111110: color_data = 8'b11111111;
		20'b00000010110000111111: color_data = 8'b11111111;
		20'b00000010110001000100: color_data = 8'b11111111;
		20'b00000010110001000101: color_data = 8'b11111111;
		20'b00000010110001001011: color_data = 8'b11111111;
		20'b00000010110001001100: color_data = 8'b11111111;
		20'b00000010110001001101: color_data = 8'b11111111;
		20'b00000010110001001110: color_data = 8'b11111111;
		20'b00000010110001001111: color_data = 8'b11111111;
		20'b00000011000000010010: color_data = 8'b11111111;
		20'b00000011000000010011: color_data = 8'b11111111;
		20'b00000011000000011011: color_data = 8'b11111111;
		20'b00000011000000011111: color_data = 8'b11111111;
		20'b00000011000000100000: color_data = 8'b11111111;
		20'b00000011000000100001: color_data = 8'b11111111;
		20'b00000011000000100010: color_data = 8'b11111111;
		20'b00000011000000100011: color_data = 8'b11111111;
		20'b00000011000000100100: color_data = 8'b11111111;
		20'b00000011000000100101: color_data = 8'b11111111;
		20'b00000011000000101001: color_data = 8'b11111111;
		20'b00000011000000101010: color_data = 8'b11111111;
		20'b00000011000000101011: color_data = 8'b11111111;
		20'b00000011000000101100: color_data = 8'b11111111;
		20'b00000011000000101101: color_data = 8'b11111111;
		20'b00000011000000101110: color_data = 8'b11111111;
		20'b00000011000000110011: color_data = 8'b11111111;
		20'b00000011000000110100: color_data = 8'b11111111;
		20'b00000011000000111010: color_data = 8'b11111111;
		20'b00000011000000111011: color_data = 8'b11111111;
		20'b00000011000000111110: color_data = 8'b11111111;
		20'b00000011000000111111: color_data = 8'b11111111;
		20'b00000011000001000100: color_data = 8'b11111111;
		20'b00000011000001000101: color_data = 8'b11111111;
		20'b00000011000001001100: color_data = 8'b11111111;
		20'b00000011000001001101: color_data = 8'b11111111;
		20'b00000011000001001110: color_data = 8'b11111111;
		20'b00000011000001001111: color_data = 8'b11111111;
		20'b00000011000001010000: color_data = 8'b11111111;
		20'b00000011000001010001: color_data = 8'b11111111;
		20'b00000011010000010011: color_data = 8'b11111111;
		20'b00000011010000010100: color_data = 8'b11111111;
		20'b00000011010000010101: color_data = 8'b11111111;
		20'b00000011010000011010: color_data = 8'b11111111;
		20'b00000011010000011011: color_data = 8'b11111111;
		20'b00000011010000011111: color_data = 8'b11111111;
		20'b00000011010000100000: color_data = 8'b11111111;
		20'b00000011010000100010: color_data = 8'b11111111;
		20'b00000011010000100011: color_data = 8'b11111111;
		20'b00000011010000100100: color_data = 8'b11111111;
		20'b00000011010000101001: color_data = 8'b11111111;
		20'b00000011010000101010: color_data = 8'b11111111;
		20'b00000011010000110011: color_data = 8'b11111111;
		20'b00000011010000110100: color_data = 8'b11111111;
		20'b00000011010000111001: color_data = 8'b11111111;
		20'b00000011010000111010: color_data = 8'b11111111;
		20'b00000011010000111011: color_data = 8'b11111111;
		20'b00000011010000111110: color_data = 8'b11111111;
		20'b00000011010000111111: color_data = 8'b11111111;
		20'b00000011010001000100: color_data = 8'b11111111;
		20'b00000011010001000101: color_data = 8'b11111111;
		20'b00000011010001001011: color_data = 8'b11111111;
		20'b00000011010001010000: color_data = 8'b11111111;
		20'b00000011010001010001: color_data = 8'b11111111;
		20'b00000011100000010011: color_data = 8'b11111111;
		20'b00000011100000010100: color_data = 8'b11111111;
		20'b00000011100000010101: color_data = 8'b11111111;
		20'b00000011100000010110: color_data = 8'b11111111;
		20'b00000011100000010111: color_data = 8'b11111111;
		20'b00000011100000011000: color_data = 8'b11111111;
		20'b00000011100000011001: color_data = 8'b11111111;
		20'b00000011100000011010: color_data = 8'b11111111;
		20'b00000011100000011011: color_data = 8'b11111111;
		20'b00000011100000011100: color_data = 8'b11111111;
		20'b00000011100000011111: color_data = 8'b11111111;
		20'b00000011100000100000: color_data = 8'b11111111;
		20'b00000011100000100100: color_data = 8'b11111111;
		20'b00000011100000100101: color_data = 8'b11111111;
		20'b00000011100000101001: color_data = 8'b11111111;
		20'b00000011100000101010: color_data = 8'b11111111;
		20'b00000011100000101011: color_data = 8'b11111111;
		20'b00000011100000101100: color_data = 8'b11111111;
		20'b00000011100000101101: color_data = 8'b11111111;
		20'b00000011100000101110: color_data = 8'b11111111;
		20'b00000011100000101111: color_data = 8'b11111111;
		20'b00000011100000110000: color_data = 8'b11111111;
		20'b00000011100000110011: color_data = 8'b11111111;
		20'b00000011100000110100: color_data = 8'b11111111;
		20'b00000011100000110101: color_data = 8'b11111111;
		20'b00000011100000110110: color_data = 8'b11111111;
		20'b00000011100000110111: color_data = 8'b11111111;
		20'b00000011100000111000: color_data = 8'b11111111;
		20'b00000011100000111001: color_data = 8'b11111111;
		20'b00000011100000111010: color_data = 8'b11111111;
		20'b00000011100000111110: color_data = 8'b11111111;
		20'b00000011100000111111: color_data = 8'b11111111;
		20'b00000011100001000100: color_data = 8'b11111111;
		20'b00000011100001000101: color_data = 8'b11111111;
		20'b00000011100001001011: color_data = 8'b11111111;
		20'b00000011100001001100: color_data = 8'b11111111;
		20'b00000011100001001101: color_data = 8'b11111111;
		20'b00000011100001001110: color_data = 8'b11111111;
		20'b00000011100001001111: color_data = 8'b11111111;
		20'b00000011100001010000: color_data = 8'b11111111;
		20'b00000011100001010001: color_data = 8'b11111111;
		20'b00000011110000010101: color_data = 8'b11111111;
		20'b00000011110000010110: color_data = 8'b11111111;
		20'b00000011110000010111: color_data = 8'b11111111;
		20'b00000011110000011000: color_data = 8'b11111111;
		20'b00000011110000011001: color_data = 8'b11111111;
		20'b00000011110000011111: color_data = 8'b11111111;
		20'b00000011110000100000: color_data = 8'b11111111;
		20'b00000011110000100100: color_data = 8'b11111111;
		20'b00000011110000100101: color_data = 8'b11111111;
		20'b00000011110000100110: color_data = 8'b11111111;
		20'b00000011110000100111: color_data = 8'b11111111;
		20'b00000011110000101001: color_data = 8'b11111111;
		20'b00000011110000101010: color_data = 8'b11111111;
		20'b00000011110000101011: color_data = 8'b11111111;
		20'b00000011110000101100: color_data = 8'b11111111;
		20'b00000011110000101101: color_data = 8'b11111111;
		20'b00000011110000101110: color_data = 8'b11111111;
		20'b00000011110000101111: color_data = 8'b11111111;
		20'b00000011110000110000: color_data = 8'b11111111;
		20'b00000011110000110011: color_data = 8'b11111111;
		20'b00000011110000110100: color_data = 8'b11111111;
		20'b00000011110000110101: color_data = 8'b11111111;
		20'b00000011110000110110: color_data = 8'b11111111;
		20'b00000011110000110111: color_data = 8'b11111111;
		20'b00000011110000111000: color_data = 8'b11111111;
		20'b00000011110000111001: color_data = 8'b11111111;
		20'b00000011110000111110: color_data = 8'b11111111;
		20'b00000011110000111111: color_data = 8'b11111111;
		20'b00000011110001000100: color_data = 8'b11111111;
		20'b00000011110001000101: color_data = 8'b11111111;
		20'b00000011110001001100: color_data = 8'b11111111;
		20'b00000011110001001101: color_data = 8'b11111111;
		20'b00000011110001001110: color_data = 8'b11111111;
		20'b00000011110001001111: color_data = 8'b11111111;
		20'b00000011110001010000: color_data = 8'b11111111;
		default: color_data = 8'b00000000;
	endcase
endmodule