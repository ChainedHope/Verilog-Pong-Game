module game_over_rom
	(
		input wire clk,
		input wire [9:0] xpos,
		input wire [9:0] ypos,
		output reg [2:0] red,
		output reg [2:0] green,
		output reg [1:0] blue
	);

	(* rom_style = "block" *)


	reg [9:0] ypos_reg;
	reg [9:0] xpos_reg;

	always @(posedge clk)
		begin
		ypos_reg <= ypos;
		xpos_reg <= xpos;
		end

	always @*
	case ({xpos_reg, ypos_reg})
		20'b00000001000000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001000000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001010000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001100000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000001110000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010010000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010100000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000010110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011100000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000011110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000100110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101000001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101100001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000010000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000101110001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110000000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110010000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000110110000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111000000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111010000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111100001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000111100001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000111110000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00000111110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000010001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000010001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000010001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000010000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110000111100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001001010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001100001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001001110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010000001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001010000001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001010000001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001010000001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001010010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010010001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001010010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001010100000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010100001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001010110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010110001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001011110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001011110001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001011110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000001010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100010001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001100010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001100100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001100100001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001100100001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100110000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001100110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001101000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001101110001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001101110001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001110000000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001110000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001110010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001110100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001110100001010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001110100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001110100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001110110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001110110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001111000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001111100001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001111100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000000000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000000001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000010000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000010001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010000010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010000100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001000001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001000001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010100001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b10; end
		20'b00010010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010110001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011000001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010011000001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011010001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010011010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010011110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010011110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100000001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100000001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010100010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010100100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010100110001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010100110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010101100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010101100001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010101110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010101110001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010101110001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010101110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110010001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010110010001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110010001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110100001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010001010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000000001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000010000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000100001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000100001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000110001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001000001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011001000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011001100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011001110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011001110001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001110001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010010001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010010001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010100001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011010110001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011010110001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010110001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011010110001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011011000000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011011000001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011011100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100000000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100010000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100010000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100100001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011100100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101000001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011101010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011101010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101100001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101110001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110000001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011110000001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011110100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111000001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111000001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011111010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011111100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011111110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000000001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000000001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000000001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000000001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000000001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000000001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100000110001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110001010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000110001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100001000000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001000001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001010000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001110001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100010010000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100010100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100010110000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100010110001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100010110001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100010110001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011000000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100011100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100011110000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100011110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100000000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100010000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100100110000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101010000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100101110000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110000000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110010000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100110110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00100111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101000110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101001110000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001110000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011100000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011100000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101011110000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011110000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101100110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101101110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101110110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110000110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110001110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110010110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110100110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000001111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101100000111100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000001111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000010000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00110101110000111101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000111100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110000000111101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011100000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011110000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100010000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111100110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111101110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110000000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110100000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111110110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010001001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b00111111110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000010000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000100000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000000110000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001000000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001010000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001100001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000001100001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000001110000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000010010001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000010010001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000010010001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000010010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000010010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010100000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000010000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000011010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011100001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011100001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000011110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000100000001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000100000001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000100000001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000100010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100010001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000100010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000100100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000100110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000100110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000100110001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000100110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000101110001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000101110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000001010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110010001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000110100000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000110100001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000110100001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111000000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111010000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111110000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111110000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111110000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111110000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111110000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111110000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111110001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000111110001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000111110001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000111110001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000000001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001000000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001000010001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001000100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001000100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001000110000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001000000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001001000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001010000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001100000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001001100001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001001100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001010000001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001010010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001010100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001010100001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001010100001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001010100001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001010100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001010110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001010110001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001010110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001011000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001011000001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001011010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001011010001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001011100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001011110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001100010001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001100010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100001010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001100110001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001100110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001101000000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001101000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001101000001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001101110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110000001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110000001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110010000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110110001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110110001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110110001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001111110000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01001111110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000000001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010000000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010000010000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000100001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010000100001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01010000100001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01010000100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010000110000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010000110001010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01010000110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01010001000000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001000001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010001000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010001000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010001010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01010001010001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01010001010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010001110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010010000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01010010010001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01010010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100001010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010010100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010010110001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01010010110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01010011000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010011000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01010011000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01010011000001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011010000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011100000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010011110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010011110000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010011110000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010100000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010100000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010100000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010100000000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010100000001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010100000001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010100010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010100010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010100010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010100100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010100100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010100110000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010100110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010100110001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010100110001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010100110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010100110001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010100110001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010100110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010101010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010101010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010101010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010101010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010101010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01010101110000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010101110000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010110000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110000000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110000000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110000001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010110000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010110010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110100001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01010110100001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010110100001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010110100001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010110100001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010110100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010110100001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01010110100001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01010110110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010110110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010110110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010110110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010110110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010110110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010110110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010110110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010110110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010111010001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b10; end
		20'b01010111010001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010001010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01010111010001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01010111100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01010111110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000000001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011000000001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011000000001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011000000001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011000000001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011000000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011000010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011000100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011000100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011000100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011000100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011000110001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011001000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011001010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001010001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011001010001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011001100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011001110001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011001110001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011010000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011010000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011010000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011010000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011010000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011010000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010100001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011010100001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011010100001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011010100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011010100001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011010100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011011000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011011010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011011100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011011110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011011110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011011110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011100000001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011100000001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b10; end
		20'b01011100010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100010001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011100010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011100010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011100010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011100010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011100010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011100010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011100110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100110001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011100110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100110001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011100110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011100110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101110001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011101110001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011101110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011101110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011110000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011110000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011110000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011110000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011110010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010001010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011110010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011110010001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01011110100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011110110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111100001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011111100001010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01011111100001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01011111100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011111100001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01011111110000001111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000010000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110000111100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01011111110001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01011111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011111110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011111110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01011111110001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011111110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01011111110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000000000001111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000010000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000111100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000000111101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000000001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100000000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000000001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100000010000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000111100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010000111101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100000110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001000001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100001000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001000001010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01100001000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100001000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001000001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01100001000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001010001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100001010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100001010001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100001100001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100001100001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100001100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100001100001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100001110001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01100001110001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01100001110001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01100001110001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01100010000000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010000000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100010000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100010010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010010000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010010000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010010001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01100010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100010010001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100010010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010010001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01100010100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010100001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100010100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011100001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100011100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011100001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01100011100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100011110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100011110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100011110001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100011110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100011110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100000001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100100000001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100100010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100010001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01100100010001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01100100100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100100001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100100100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100100100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100100100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100100100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100100100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100100100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000101011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000101110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000110001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100100110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100100110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101000001010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101000001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100101000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100101010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100101010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101010001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01100101100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101100001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01100101110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100101110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100110000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100110000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110000001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100110000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110010001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110010001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100110010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100110010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100110100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100110100001010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01100110100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100110110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100110110001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01100110110001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01100111000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100111000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100111000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100111000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100111000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100111000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01100111000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111100001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100111100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01100111100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01100111110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01100111110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101000000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100000101111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101000100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101000100001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101000100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101000110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101000110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000000110010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000001010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101001000001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101001000001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101001010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001010001010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01101001010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01101001100000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101001100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001100001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101001100001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101001100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101001100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101001100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101001100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101001100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001110000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110000111011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101001110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101001110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010000000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000101010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010000001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010000001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010010000010001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000101011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000101100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010100000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000101001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000101100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000101101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010100001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010110000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000101101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000101110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101010110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101010110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011000000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000101111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000110000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101011000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011010000010010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000101000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000110000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000110001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101011100000010011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000110010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000110011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100001010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101011100001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101011100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101011110000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000100111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000110100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101011110001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01101011110001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01101100000000010100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000100110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000110101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000110110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101100000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101100000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101100000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101100000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101100000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101100000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100010000010101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000010110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000100101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000110111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100010001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100100000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000010111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000011000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000100011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000100100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000110111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000111000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100001010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101100100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01101100100001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101100110000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000011001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000011010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000011011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000011100: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000011101: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000011110: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000011111: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000100000: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000100001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000100010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000111001: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110001010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101100110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101100110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01101101000000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000000011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000000011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000000011101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000000011110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000000011111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000000100000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000000111010: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101101000001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101000001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01101101010000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101101010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101101010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01101101100000111011: begin red <= 3'b111; green <= 3'b000; blue <= 2'b00; end
		20'b01101101100001010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01101101100001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01101101100001010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01101101100001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01101101100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101101100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101101110001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101101110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101110000001010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101110000001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101110000001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101110000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101110000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101110000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101110000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01101110000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01101110010001010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01101110010001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		default: begin red <= 3'b000; green <= 3'b000; blue <= 2'b00; end
	endcase
endmodule