module pong_menu_rom
	(
		input wire clk,
		input wire [9:0] row,
		input wire [9:0] col,
		output reg [7:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [9:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})








		20'b00000010000000010001: color_data = 8'b11111111;
		20'b00000010000000010010: color_data = 8'b11111111;
		20'b00000010000000010011: color_data = 8'b11111111;
		20'b00000010000000010100: color_data = 8'b11111111;
		20'b00000010000000010101: color_data = 8'b11111111;
		20'b00000010000000010110: color_data = 8'b11111111;
		20'b00000010000000010111: color_data = 8'b11111111;
		20'b00000010000000011000: color_data = 8'b11111111;
		20'b00000010000000011111: color_data = 8'b11111111;
		20'b00000010000000100000: color_data = 8'b11111111;
		20'b00000010000000100001: color_data = 8'b11111111;
		20'b00000010000000100010: color_data = 8'b11111111;
		20'b00000010000000100011: color_data = 8'b11111111;
		20'b00000010000000101001: color_data = 8'b11111111;
		20'b00000010000000101010: color_data = 8'b11111111;
		20'b00000010000000101011: color_data = 8'b11111111;
		20'b00000010000000110001: color_data = 8'b11111111;
		20'b00000010000000110010: color_data = 8'b11111111;
		20'b00000010000000110011: color_data = 8'b11111111;
		20'b00000010000000111001: color_data = 8'b11111111;
		20'b00000010000000111010: color_data = 8'b11111111;
		20'b00000010000000111011: color_data = 8'b11111111;
		20'b00000010000000111100: color_data = 8'b11111111;
		20'b00000010000000111101: color_data = 8'b11111111;

		20'b00000010010000010001: color_data = 8'b11111111;
		20'b00000010010000010010: color_data = 8'b11111111;
		20'b00000010010000010011: color_data = 8'b11111111;
		20'b00000010010000010100: color_data = 8'b11111111;
		20'b00000010010000010101: color_data = 8'b11111111;
		20'b00000010010000010110: color_data = 8'b11111111;
		20'b00000010010000010111: color_data = 8'b11111111;
		20'b00000010010000011000: color_data = 8'b11111111;
		20'b00000010010000011001: color_data = 8'b11111111;
		20'b00000010010000011101: color_data = 8'b11111111;
		20'b00000010010000011110: color_data = 8'b11111111;
		20'b00000010010000011111: color_data = 8'b11111111;
		20'b00000010010000100000: color_data = 8'b11111111;
		20'b00000010010000100001: color_data = 8'b11111111;
		20'b00000010010000100010: color_data = 8'b11111111;
		20'b00000010010000100011: color_data = 8'b11111111;
		20'b00000010010000100100: color_data = 8'b11111111;
		20'b00000010010000100101: color_data = 8'b11111111;
		20'b00000010010000101001: color_data = 8'b11111111;
		20'b00000010010000101010: color_data = 8'b11111111;
		20'b00000010010000101011: color_data = 8'b11111111;
		20'b00000010010000101100: color_data = 8'b11111111;
		20'b00000010010000110010: color_data = 8'b11111111;
		20'b00000010010000110011: color_data = 8'b11111111;
		20'b00000010010000110111: color_data = 8'b11111111;
		20'b00000010010000111000: color_data = 8'b11111111;
		20'b00000010010000111001: color_data = 8'b11111111;
		20'b00000010010000111010: color_data = 8'b11111111;
		20'b00000010010000111011: color_data = 8'b11111111;
		20'b00000010010000111100: color_data = 8'b11111111;
		20'b00000010010000111101: color_data = 8'b11111111;
		20'b00000010010000111110: color_data = 8'b11111111;
		20'b00000010010000111111: color_data = 8'b11111111;

		20'b00000010100000010001: color_data = 8'b11111111;
		20'b00000010100000010010: color_data = 8'b11111111;
		20'b00000010100000010011: color_data = 8'b11111111;
		20'b00000010100000011000: color_data = 8'b11111111;
		20'b00000010100000011001: color_data = 8'b11111111;
		20'b00000010100000011010: color_data = 8'b11111111;
		20'b00000010100000011100: color_data = 8'b11111111;
		20'b00000010100000011101: color_data = 8'b11111111;
		20'b00000010100000011110: color_data = 8'b11111111;
		20'b00000010100000011111: color_data = 8'b11111111;
		20'b00000010100000100011: color_data = 8'b11111111;
		20'b00000010100000100100: color_data = 8'b11111111;
		20'b00000010100000100101: color_data = 8'b11111111;
		20'b00000010100000100110: color_data = 8'b11111111;
		20'b00000010100000101001: color_data = 8'b11111111;
		20'b00000010100000101010: color_data = 8'b11111111;
		20'b00000010100000101011: color_data = 8'b11111111;
		20'b00000010100000101100: color_data = 8'b11111111;
		20'b00000010100000101101: color_data = 8'b11111111;
		20'b00000010100000110010: color_data = 8'b11111111;
		20'b00000010100000110011: color_data = 8'b11111111;
		20'b00000010100000110110: color_data = 8'b11111111;
		20'b00000010100000110111: color_data = 8'b11111111;
		20'b00000010100000111000: color_data = 8'b11111111;
		20'b00000010100000111001: color_data = 8'b11111111;
		20'b00000010100000111110: color_data = 8'b11111111;
		20'b00000010100000111111: color_data = 8'b11111111;

		20'b00000010110000010001: color_data = 8'b11111111;
		20'b00000010110000010010: color_data = 8'b11111111;
		20'b00000010110000010011: color_data = 8'b11111111;
		20'b00000010110000011000: color_data = 8'b11111111;
		20'b00000010110000011001: color_data = 8'b11111111;
		20'b00000010110000011010: color_data = 8'b11111111;
		20'b00000010110000011100: color_data = 8'b11111111;
		20'b00000010110000011101: color_data = 8'b11111111;
		20'b00000010110000100101: color_data = 8'b11111111;
		20'b00000010110000100110: color_data = 8'b11111111;
		20'b00000010110000101001: color_data = 8'b11111111;
		20'b00000010110000101010: color_data = 8'b11111111;
		20'b00000010110000101011: color_data = 8'b11111111;
		20'b00000010110000101100: color_data = 8'b11111111;
		20'b00000010110000101101: color_data = 8'b11111111;
		20'b00000010110000101110: color_data = 8'b11111111;
		20'b00000010110000110010: color_data = 8'b11111111;
		20'b00000010110000110011: color_data = 8'b11111111;
		20'b00000010110000110110: color_data = 8'b11111111;
		20'b00000010110000110111: color_data = 8'b11111111;

		20'b00000011000000010001: color_data = 8'b11111111;
		20'b00000011000000010010: color_data = 8'b11111111;
		20'b00000011000000010011: color_data = 8'b11111111;
		20'b00000011000000010100: color_data = 8'b11111111;
		20'b00000011000000010101: color_data = 8'b11111111;
		20'b00000011000000010110: color_data = 8'b11111111;
		20'b00000011000000010111: color_data = 8'b11111111;
		20'b00000011000000011000: color_data = 8'b11111111;
		20'b00000011000000011001: color_data = 8'b11111111;
		20'b00000011000000011100: color_data = 8'b11111111;
		20'b00000011000000011101: color_data = 8'b11111111;
		20'b00000011000000100101: color_data = 8'b11111111;
		20'b00000011000000100110: color_data = 8'b11111111;
		20'b00000011000000101001: color_data = 8'b11111111;
		20'b00000011000000101010: color_data = 8'b11111111;
		20'b00000011000000101101: color_data = 8'b11111111;
		20'b00000011000000101110: color_data = 8'b11111111;
		20'b00000011000000101111: color_data = 8'b11111111;
		20'b00000011000000110010: color_data = 8'b11111111;
		20'b00000011000000110011: color_data = 8'b11111111;
		20'b00000011000000110110: color_data = 8'b11111111;
		20'b00000011000000110111: color_data = 8'b11111111;

		20'b00000011010000010001: color_data = 8'b11111111;
		20'b00000011010000010010: color_data = 8'b11111111;
		20'b00000011010000010011: color_data = 8'b11111111;
		20'b00000011010000010100: color_data = 8'b11111111;
		20'b00000011010000010101: color_data = 8'b11111111;
		20'b00000011010000010110: color_data = 8'b11111111;
		20'b00000011010000010111: color_data = 8'b11111111;
		20'b00000011010000011000: color_data = 8'b11111111;
		20'b00000011010000011100: color_data = 8'b11111111;
		20'b00000011010000011101: color_data = 8'b11111111;
		20'b00000011010000100101: color_data = 8'b11111111;
		20'b00000011010000100110: color_data = 8'b11111111;
		20'b00000011010000101001: color_data = 8'b11111111;
		20'b00000011010000101010: color_data = 8'b11111111;
		20'b00000011010000101110: color_data = 8'b11111111;
		20'b00000011010000101111: color_data = 8'b11111111;
		20'b00000011010000110000: color_data = 8'b11111111;
		20'b00000011010000110010: color_data = 8'b11111111;
		20'b00000011010000110011: color_data = 8'b11111111;
		20'b00000011010000110110: color_data = 8'b11111111;
		20'b00000011010000110111: color_data = 8'b11111111;
		20'b00000011010000111011: color_data = 8'b11111111;
		20'b00000011010000111100: color_data = 8'b11111111;
		20'b00000011010000111101: color_data = 8'b11111111;
		20'b00000011010000111110: color_data = 8'b11111111;
		20'b00000011010000111111: color_data = 8'b11111111;
		20'b00000011010001000000: color_data = 8'b11111111;

		20'b00000011100000010001: color_data = 8'b11111111;
		20'b00000011100000010010: color_data = 8'b11111111;
		20'b00000011100000010011: color_data = 8'b11111111;
		20'b00000011100000011100: color_data = 8'b11111111;
		20'b00000011100000011101: color_data = 8'b11111111;
		20'b00000011100000100101: color_data = 8'b11111111;
		20'b00000011100000100110: color_data = 8'b11111111;
		20'b00000011100000101001: color_data = 8'b11111111;
		20'b00000011100000101010: color_data = 8'b11111111;
		20'b00000011100000101111: color_data = 8'b11111111;
		20'b00000011100000110000: color_data = 8'b11111111;
		20'b00000011100000110001: color_data = 8'b11111111;
		20'b00000011100000110010: color_data = 8'b11111111;
		20'b00000011100000110011: color_data = 8'b11111111;
		20'b00000011100000110110: color_data = 8'b11111111;
		20'b00000011100000110111: color_data = 8'b11111111;
		20'b00000011100000111011: color_data = 8'b11111111;
		20'b00000011100000111100: color_data = 8'b11111111;
		20'b00000011100000111101: color_data = 8'b11111111;
		20'b00000011100000111110: color_data = 8'b11111111;
		20'b00000011100000111111: color_data = 8'b11111111;
		20'b00000011100001000000: color_data = 8'b11111111;

		20'b00000011110000010001: color_data = 8'b11111111;
		20'b00000011110000010010: color_data = 8'b11111111;
		20'b00000011110000010011: color_data = 8'b11111111;
		20'b00000011110000011100: color_data = 8'b11111111;
		20'b00000011110000011101: color_data = 8'b11111111;
		20'b00000011110000011110: color_data = 8'b11111111;
		20'b00000011110000011111: color_data = 8'b11111111;
		20'b00000011110000100011: color_data = 8'b11111111;
		20'b00000011110000100100: color_data = 8'b11111111;
		20'b00000011110000100101: color_data = 8'b11111111;
		20'b00000011110000100110: color_data = 8'b11111111;
		20'b00000011110000101001: color_data = 8'b11111111;
		20'b00000011110000101010: color_data = 8'b11111111;
		20'b00000011110000110000: color_data = 8'b11111111;
		20'b00000011110000110001: color_data = 8'b11111111;
		20'b00000011110000110010: color_data = 8'b11111111;
		20'b00000011110000110011: color_data = 8'b11111111;
		20'b00000011110000110110: color_data = 8'b11111111;
		20'b00000011110000110111: color_data = 8'b11111111;
		20'b00000011110000111000: color_data = 8'b11111111;
		20'b00000011110000111001: color_data = 8'b11111111;
		20'b00000011110000111111: color_data = 8'b11111111;
		20'b00000011110001000000: color_data = 8'b11111111;

		20'b00000100000000010001: color_data = 8'b11111111;
		20'b00000100000000010010: color_data = 8'b11111111;
		20'b00000100000000010011: color_data = 8'b11111111;
		20'b00000100000000011101: color_data = 8'b11111111;
		20'b00000100000000011110: color_data = 8'b11111111;
		20'b00000100000000011111: color_data = 8'b11111111;
		20'b00000100000000100000: color_data = 8'b11111111;
		20'b00000100000000100001: color_data = 8'b11111111;
		20'b00000100000000100010: color_data = 8'b11111111;
		20'b00000100000000100011: color_data = 8'b11111111;
		20'b00000100000000100100: color_data = 8'b11111111;
		20'b00000100000000100101: color_data = 8'b11111111;
		20'b00000100000000101001: color_data = 8'b11111111;
		20'b00000100000000101010: color_data = 8'b11111111;
		20'b00000100000000110001: color_data = 8'b11111111;
		20'b00000100000000110010: color_data = 8'b11111111;
		20'b00000100000000110011: color_data = 8'b11111111;
		20'b00000100000000110111: color_data = 8'b11111111;
		20'b00000100000000111000: color_data = 8'b11111111;
		20'b00000100000000111001: color_data = 8'b11111111;
		20'b00000100000000111010: color_data = 8'b11111111;
		20'b00000100000000111011: color_data = 8'b11111111;
		20'b00000100000000111100: color_data = 8'b11111111;
		20'b00000100000000111101: color_data = 8'b11111111;
		20'b00000100000000111110: color_data = 8'b11111111;
		20'b00000100000000111111: color_data = 8'b11111111;

		20'b00000100010000010001: color_data = 8'b11111111;
		20'b00000100010000010010: color_data = 8'b11111111;
		20'b00000100010000010011: color_data = 8'b11111111;
		20'b00000100010000011111: color_data = 8'b11111111;
		20'b00000100010000100000: color_data = 8'b11111111;
		20'b00000100010000100001: color_data = 8'b11111111;
		20'b00000100010000100010: color_data = 8'b11111111;
		20'b00000100010000100011: color_data = 8'b11111111;
		20'b00000100010000101001: color_data = 8'b11111111;
		20'b00000100010000101010: color_data = 8'b11111111;
		20'b00000100010000101011: color_data = 8'b11111111;
		20'b00000100010000110001: color_data = 8'b11111111;
		20'b00000100010000110010: color_data = 8'b11111111;
		20'b00000100010000110011: color_data = 8'b11111111;
		20'b00000100010000111001: color_data = 8'b11111111;
		20'b00000100010000111010: color_data = 8'b11111111;
		20'b00000100010000111011: color_data = 8'b11111111;
		20'b00000100010000111100: color_data = 8'b11111111;
		20'b00000100010000111101: color_data = 8'b11111111;






		default: color_data = 8'b00000000;
	endcase
endmodule