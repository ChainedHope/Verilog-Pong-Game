module credits_rom
	(
		input wire clk,
		input wire [9:0] xpos,
		input wire [9:0] ypos,
		output reg [2:0] red,
		output reg [2:0] green,
		output reg [1:0] blue
	);

	(* rom_style = "block" *)


	reg [9:0] ypos_reg;
	reg [9:0] xpos_reg;

	always @(posedge clk)
		begin
		ypos_reg <= ypos;
		xpos_reg <= xpos;
		end

	always @*
	case ({xpos_reg, ypos_reg})
		20'b00000000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011010000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011010000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000011010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000011010000111001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000011010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011100000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011100000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011100000110111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000011100000111000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000011100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000110101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000011110000110110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000011110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000100000000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000100000000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000100000000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000100000000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000100000000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000100000000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000100000000011010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100000000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000100000000110100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000100000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100000000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100000000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000110001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010000110010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000100010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000100100000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000100100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000100110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110000110101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000100110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000101000000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000101000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000110001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000101000000110010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000101000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000101010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000101010000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000101010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101010000111001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000101010000111010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100000010001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000101100000010010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000101100000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000101100000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000101100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000101100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000101100000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000101100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000101110000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000101110000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000101110000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00000101110000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000101110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110010000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000110010000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000110100000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000110100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00000110100000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000110100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000110110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000111000000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00000111000000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111000000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111000000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111000000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111000000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000101010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000010011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000111100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000111100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000111100000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00000111100000011010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111110000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00000111110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00000111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00000111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000000000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000000000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000000000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001000000000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001000000000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001000010000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001000010000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000010000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001000010000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001000010000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001000100000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000100000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000100000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000100000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000100000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000100000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001000100000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001000100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000100000101001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001000100000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000100000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000110000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001000110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001000110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001001000000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001001000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001001010000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001001010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001001010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001001010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001001100000010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001001100000010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001001100000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001001100000011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001001100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001001110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000011010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001010000000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001010000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010010000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001010110000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010110000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010110000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001010110000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001010110000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001011000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011000000010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001011000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001011000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011000000011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001011000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011000000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001011000000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001011000000110011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001011010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001011010000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001011010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001011010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010000110100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001011010000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001011100000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001011100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001011100000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001011100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011100000110101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001011100000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001011110000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001011110000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000100011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000000100100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001100000000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001100000000100110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001100000000100111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001100000000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001100000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100000000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001100000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100000000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100010000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001100010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100010000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100100000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100100000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100100000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100100000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100100000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100100000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001100100000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100100000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100000111010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001100110000010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001100110000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001100110000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001100110000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001100110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100110000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001100110000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001100110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001101000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001101000000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001101000000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001101000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001101000000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001101000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001101010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001101010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001101010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001101010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001101010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001101100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001101100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100000111001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001101100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001101110000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001101110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001101110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001101110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000110111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001101110000111000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001101110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000110101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001110000000110110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001110000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110000000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000110011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010000110100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001110010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001110010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001110100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001110100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001110100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001110110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001110110000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001110110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110000110111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001110110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001111000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001111000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111000000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111000000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00001111000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111000000111010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111010000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111010000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001111010000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001111010000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111010000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001111100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111100000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001111100000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001111100000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001111100000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001111100000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00001111100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00001111110000011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00001111110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00001111110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00001111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00001111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010000000000010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010000000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010000000000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010000000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000000000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010000000000110011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010000000000111010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010000010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010000010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000010000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010000110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010000110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010000110000110110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010000110000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001000000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010001000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010001000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001000000110111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010001010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001010000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010001010000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001010000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001100000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010001100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001100000111001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001100001010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001100001011100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010001110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001110000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010001110000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010001110000110011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010001110000110100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001110000110101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001110000110110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010001110000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010001110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110000111010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010001110001010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010001110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010010000000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010000000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010000000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010000000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010000000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010000000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010000000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010010000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010010000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010010000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010010000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010010000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010010000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010010001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010001011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010010001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010100000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010100000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010100000100110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010100000100111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010100000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010100000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010100000101010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010010100000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010110000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010010110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010010110000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010110000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010010110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010010110000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010110000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000000011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010011000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011000000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011000000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011000000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010011010001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010011010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010011100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011100000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010011100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011100000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011100000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011100000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011100001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011110000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010011110000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010011110000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010011110000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011110000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010011110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010011110001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011110001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011110001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010011110001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100000001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010100000001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010100000001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010100000001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010100000001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010100000001011011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010100000001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100000110101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010100100000111000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010100100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100100001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010100110000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010100110001011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010101000000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010101000000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101000001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101000001011100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101010000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010101010000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010101010000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010101010000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101100000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010101100000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010101100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010101110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010101110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010101110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010101110001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010101110001011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010101110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010110000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110000001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110000001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110010001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010110010001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010110010001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010110010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010110010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010110010001011011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010110010001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110110000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010110110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010110110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010110110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010110110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00010111000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111010000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111010000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111010000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111010000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111010000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111010000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00010111010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111010000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00010111100000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111100000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00010111110000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00010111110000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111110000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00010111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00010111110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000000000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000000000110011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000000000111010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011000000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011000000001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011000000001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000010000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000010000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000010000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000010001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000010001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000010001011011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000100000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000100000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000100000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000100000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000100000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100000101001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011000100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000100001011100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011000110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011000110000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011000110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011000110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011001000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011001000000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011001000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011001000000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011001000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001000000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001000000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001000000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011001010000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011001010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011001010000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011001010000011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011001010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001010000111001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001100000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011001100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011001100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011001100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100000111010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011001100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011001100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011001110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011001110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011001110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011001110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011001110001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011010000000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010000000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010000000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010000000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010000001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010000001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010000001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000010011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010010000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011010010000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011010010000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010010000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010010000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011010010000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010010000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010010001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010010001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011010010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011010010001011011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011010100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010100001011100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011010110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011011000000100001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011000000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011010000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011010000100010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000101001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100000110001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011100000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011011110000011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110000100010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011011110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110000110010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000110011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011011110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011011110001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011100000000010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100000000100001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100000001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011100000001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100000001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000010011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011100010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100010000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100010000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100010000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011100100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011100110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011101000000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011101000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011101000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011101000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101000000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011101010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101010000111001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101010000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011101100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000110001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101100000110100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011101100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011101110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011101110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110000110001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011101110000110010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011101110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011101110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011110000000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011110000000100111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011110000000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110000000110010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110000000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110000000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011110000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011110010000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110010000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00011110010000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110010001011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000100011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011110100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110100000110101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011110100000110110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110100000110111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110100000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011110110000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011110110000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011110110000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011110110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011110110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000110100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011110110000111001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011110110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011111000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011111000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111000000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111010000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111010000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111010000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111110000011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00011111110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00011111110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00011111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00011111110001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00011111110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100000000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100000000000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010000110101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000111000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000010001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000010001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000010001011011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000010001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100000100000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100000100000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100000100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000110000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100000110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100000110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100000110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100000110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001000000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001000000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100001000000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100001000000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001000001011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001010000110011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001010000110100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001010000110101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001010000110110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001010000110111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001010000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001010000111001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001010000111010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100001100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100001100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000101010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100001110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100001110001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100001110001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010000000110111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010000000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100010000000111010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010000001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010010000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010010000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010000111001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010010001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010100000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100010100000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010100000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010100000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000110101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100010110000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100010110000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100010110000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100010110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011000000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100011000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100011000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011000000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011000000110011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011000000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100011000000111001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100011000000111010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100011010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011010001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100011100000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100011100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011100001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100011110000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100011110000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100011110000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100011110001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100011110001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100011110001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100000000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100010000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100010000101010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100100010000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100100100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100100110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100100110000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100100110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100100110001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100100110001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100100110001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100101000000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100101000000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100101000000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100101000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100101000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101000001011011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100101010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100101100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101100001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100101110000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100101110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100101110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000101001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110000000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100110010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100110100000010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100110100000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110100000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110100000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110100000110011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100110100000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110100000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110000011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110110000110011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110110000111010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100110110001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100110110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100110110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100110110001011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100111000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100111000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100111000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100111000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100111000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000000110100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000111000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000111001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100111000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100111010000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100111010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111010001010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100111010001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100111010001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00100111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111100000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000111001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00100111100000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00100111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111100001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100111100001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100111100001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100111100001011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00100111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00100111110000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00100111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00100111110001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000000111001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101000000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000000001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101000010000011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101000010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000010000111010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000100001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101000100000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101000100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000110101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101000100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101000110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101000110000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000100010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000100011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000110011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101000110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101000110000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101000110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101000110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001000000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000000110100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001000000110110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101001000000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101001000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001000001011100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101001010000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101001010000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010000100010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001010000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001010000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001010000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001010000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010000110101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101001010000110110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101001010000110111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101001010000111000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001010001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101001100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000110100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101001100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001100000111001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001100001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001100001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001100001011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101001110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000100111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101001110000110011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101001110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101001110000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101001110000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101001110000111010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101001110001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101001110001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101010000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101010000000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101010000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101010000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000110101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101010000000111000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101010000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101010010000100001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101010010000100010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101010010000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000101001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101010010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101010010000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101010100000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101010100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010100001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101010100001011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000011010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000100010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101010110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101010110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101010110001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000100001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000100010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011000000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000110011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000110101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101011000000111000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101011000000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011010000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010000100001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101011010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101011010000110100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010000110110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000110111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101011010001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011010001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011010001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011100000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101011100000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101011100000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101011100000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101011100000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101011100000110100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011100000110101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100000110110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100000110111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100000111000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101011110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110000101001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101011110000110101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011110000110110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011110000110111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101011110000111000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101011110001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101011110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101100000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101100000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100000000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100000001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101100000001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100000001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101100010000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101100010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100010000111001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101100010000111010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100100000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100000111001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100000111010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100100001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100100001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100100001011011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101100100001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101100110000111001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101100110000111010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101100110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101101010000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101101010000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101101010000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101101010000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101101010000011010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101101010000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101101010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101010001011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101110000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101110000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101110000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101110000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101101110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101101110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101101110000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101110000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101110000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101110000000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110000001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101110000001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101110010000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101110010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101110100000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101110100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110100001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110110000100111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101110110000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101110110001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101110110001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101111000000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101111000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101111000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111000001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101111000001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00101111010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101111010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111010001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101111100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111100001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101111110000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111110000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101111110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00101111110000100110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00101111110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00101111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00101111110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00101111110001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00101111110001011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000000000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110000000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110000000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000000001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000010000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110000010000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110000010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110000010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000100000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110000100000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110000100001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110000100001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000100001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000100001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000010011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110000110000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110000110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000110000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110000110000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110000110000011010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000110000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000110001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000110001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110000110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110000110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001000001010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000001011011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001010000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110001010000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110001010000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110001010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110001010000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110001010000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110001010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001010000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110001010000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001010000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001010000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001010000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001010000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001010001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001010001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110001100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001100001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110001100001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110001100001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110001100001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110001100001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110001100001011011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110001110000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110001110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110001110001011100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010000000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110010000001011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110010000001011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110010000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110010010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110010100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110010100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110010110000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110010110000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110010110000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110010110000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110010110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110011000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000000101001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000001010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110011000001011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110011000001011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110011000001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110011010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110011010000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110011010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011010000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011010001011100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110011100000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110011100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110011100000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110011100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011100001010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011100001010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100001011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100001011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100001011010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011100001011011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110011110001010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110011110001010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110011110001011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110011110001011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110011110001011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110011110001011011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110011110001011100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110100000000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110100000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110100000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100010001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100100000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110100100000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110100100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100100001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100110000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110100110001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110101000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101000000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101000001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101000001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110101010000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110101010000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110101010000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110101010000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110101010000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101010001011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101100000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101100000100100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101100001010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110101100001010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110101100001011011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110101100001011100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110101110000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110000100110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110110000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110110000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110110000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110000000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110110000000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110110000000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110110010000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110110010000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110110010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100000100110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110110100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110110100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110110110000100100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110110110000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110110110000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110110110000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110111000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110111000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111000000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110111000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111010000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110111100000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110111100000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110111100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110111100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111100000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110111100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111100000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110111100000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110111100000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110111110000010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110111110000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00110111110000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00110111110000100011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00110111110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00110111110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00110111110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00110111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00110111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000000000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000000100110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111000000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111000000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111000010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000010000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111000010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111000010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000010000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111000010000100011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111000010000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000010000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111000010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111000100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111000100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111000100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111000110000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111000110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001000000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111001000000100100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111001000000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111001000000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111001000000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111001000000101001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111001010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111001100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111001100000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111001100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001100000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111001100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001100000101010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001110000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111001110000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111001110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111010000000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111010000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111010010000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111010010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010100000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010100000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111010100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010100000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111010100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111010100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010100000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111010100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111010110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111010110000101010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111011000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111011000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011000000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111011000000100111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111011000000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111011000000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011010000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111011010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011100000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111100000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111100000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100000000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111100000000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111100000000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100000000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100010000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100010000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100000010011: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111100100000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111100100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111100100000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111100100000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111100100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111100100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100100000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111100110000011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111100110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111100110000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111100110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111100110000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110000101010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101000000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101000000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111101000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101010000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111101010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101100000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111101100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101100000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111101100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101110000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111101110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111101110000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111101110000100100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101110000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101110000100110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101110000100111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101110000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101110000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111101110000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000000010001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111110000000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111110000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111110000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111110010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111110010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110100000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110100000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110100000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111110100000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111111000000010010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111111000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111111000000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111111000000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111111000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111111000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111111000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111111000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111111000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b00111111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010000010001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b00111111010000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111111010000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b00111111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111111100000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b00111111100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111111100000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111111100000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000010010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111111110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111111110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111111110000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111111110000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b00111111110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b00111111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b00111111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000000010001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000000000000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000000000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000000000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000000000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000000000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000000000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000000000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000000000000100111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000000000000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000000000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000000010000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000000010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000000010000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000000010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000010000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000100011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100000100100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000000100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000000100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000000110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000000100111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000001000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000010001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000001010000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000001010000010101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000001010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001010000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b10; end
		20'b01000001010000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001010000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000001010000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000001010000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000001010000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000001010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000001100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000001100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110000010010: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000001110000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000001110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001110000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000001110000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000001110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000010110: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000101001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000010000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010000010001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000010010000010010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000010010000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000010010000101010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010100000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010100000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000011010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011000000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011000000011001: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000011000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011000000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000011000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011000000100110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000011000000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011010000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011010000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000011010000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011010000100100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000011010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011010000100111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011100000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000011100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011100000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000011100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000011100000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000011100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011100000101000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011110000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011110000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000011110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011110000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000011110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000011110000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011110000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000011110000101001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100000000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100000000010011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100000000010111: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000100000000100011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000100000000100100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000100000000100101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000100000000100110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000100000000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100000000101010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000100010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100000010001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100100000010010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100100000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100100000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000100100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100100000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100100000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100100000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100100000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000100100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110000010001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000100110000010010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000100110000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000100110000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000000100011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000101000000101010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01000101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101010000100100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000100101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000101000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000101001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101100000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101100000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101100000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101100000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101110000100101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000101110000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000101110000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000101110000101000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000101110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000110000000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000110000000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110000000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110010000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110010000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110010000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110010000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110010000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110110000010101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110110000011000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000110110000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000110110000100011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110110000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110110000100101: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000110110000101000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01000110110000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110110000101010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111000000100011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000111000000100100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111000000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111000000100110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000100111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111000000101001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111000000101010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111010000100100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000111010000100101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111010000100110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111010000100111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111010000101000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111010000101001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111100000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000111100000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01000111100000100101: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100000100110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000111100000100111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01000111100000101000: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01000111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01000111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01000111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001000000000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001000010000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000010000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000010000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000010000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000010000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000010000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001000010000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000100000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000100000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001001000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001001010000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001100000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001010000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010000000010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001010000000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010000010100: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001010010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010010000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001010100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010100000011000: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001010110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001010110000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000000010011: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001011000000010100: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001011000000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001011000000010110: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001011000000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001011000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011000000011010: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011010000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011010000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011100000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001011100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001011100000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001011100000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001011100000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001011100000011001: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001011100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001011100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001011110000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001011110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001011110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000000011001: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001100000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010000010111: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001100010000011000: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001100010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100000010101: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001100100000010110: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001100100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100100000011010: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001100100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000010011: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110000010100: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001100110000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100110000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100110000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001100110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001100110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001100110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101000000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001101000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101010000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101010000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101010000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010000010111: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001101010000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001101100000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001101100000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001101100000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101100000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101100000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101100000011010: begin red <= 3'b000; green <= 3'b100; blue <= 2'b10; end
		20'b01001101100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001101110000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101110000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001101110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001101110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001110000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001110000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001110000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010000011001: begin red <= 3'b100; green <= 3'b000; blue <= 2'b00; end
		20'b01001110010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001110010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100000010011: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110100000011010: begin red <= 3'b000; green <= 3'b000; blue <= 2'b10; end
		20'b01001110100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001110110000010100: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000010101: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000010110: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000010111: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000011000: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000011001: begin red <= 3'b000; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001110110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001110110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000000010011: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000000010100: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000000010101: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000000010110: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000000010111: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000000011000: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010000010011: begin red <= 3'b100; green <= 3'b100; blue <= 2'b10; end
		20'b01001111010000010100: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001111010000010101: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001111010000010110: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001111010000010111: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001111010000011000: begin red <= 3'b100; green <= 3'b100; blue <= 2'b00; end
		20'b01001111010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111110000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01001111110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01001111110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010000000000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010000000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010000010000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010000010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100000011001: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010000100000011010: begin red <= 3'b110; green <= 3'b110; blue <= 2'b11; end
		20'b01010000100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010000110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010001110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010100001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010010110001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011000001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000001011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000001100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000001101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000001110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000001111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000010000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000010001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000010010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000010011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000010100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000010101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000010110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000010111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000011000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000011001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000011010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000011011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000011100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000011101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000011110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000011111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000100000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000100001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000100010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000100011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000100100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000100101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000100110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000100111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000101000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000101001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000101010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000101011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000101100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000101101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000101110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000101111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000110000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000110001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000110010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000110011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000110100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000110101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000110110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000110111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000111000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000111001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000111010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000111011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000111100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000111101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000111110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010000111111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001000000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001000001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001000010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001000011: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001000100: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001000101: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001000110: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001000111: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001001000: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001001001: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		20'b01010011010001001010: begin red <= 3'b111; green <= 3'b111; blue <= 2'b11; end
		default: begin red <= 3'b000; green <= 3'b000; blue <= 2'b00; end
	endcase
endmodule